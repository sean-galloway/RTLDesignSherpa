`timescale 1ns / 1ps

module math_multiplier_wallace_tree_csa_16 (
    input  [15:0] i_multiplier,
    input  [15:0] i_multiplicand,
    output [31:0] ow_product
);

// Partial products generation
wire w_pp_0_0 = i_multiplier[0] & i_multiplicand[0];
wire w_pp_0_1 = i_multiplier[0] & i_multiplicand[1];
wire w_pp_0_2 = i_multiplier[0] & i_multiplicand[2];
wire w_pp_0_3 = i_multiplier[0] & i_multiplicand[3];
wire w_pp_0_4 = i_multiplier[0] & i_multiplicand[4];
wire w_pp_0_5 = i_multiplier[0] & i_multiplicand[5];
wire w_pp_0_6 = i_multiplier[0] & i_multiplicand[6];
wire w_pp_0_7 = i_multiplier[0] & i_multiplicand[7];
wire w_pp_0_8 = i_multiplier[0] & i_multiplicand[8];
wire w_pp_0_9 = i_multiplier[0] & i_multiplicand[9];
wire w_pp_0_10 = i_multiplier[0] & i_multiplicand[10];
wire w_pp_0_11 = i_multiplier[0] & i_multiplicand[11];
wire w_pp_0_12 = i_multiplier[0] & i_multiplicand[12];
wire w_pp_0_13 = i_multiplier[0] & i_multiplicand[13];
wire w_pp_0_14 = i_multiplier[0] & i_multiplicand[14];
wire w_pp_0_15 = i_multiplier[0] & i_multiplicand[15];
wire w_pp_1_0 = i_multiplier[1] & i_multiplicand[0];
wire w_pp_1_1 = i_multiplier[1] & i_multiplicand[1];
wire w_pp_1_2 = i_multiplier[1] & i_multiplicand[2];
wire w_pp_1_3 = i_multiplier[1] & i_multiplicand[3];
wire w_pp_1_4 = i_multiplier[1] & i_multiplicand[4];
wire w_pp_1_5 = i_multiplier[1] & i_multiplicand[5];
wire w_pp_1_6 = i_multiplier[1] & i_multiplicand[6];
wire w_pp_1_7 = i_multiplier[1] & i_multiplicand[7];
wire w_pp_1_8 = i_multiplier[1] & i_multiplicand[8];
wire w_pp_1_9 = i_multiplier[1] & i_multiplicand[9];
wire w_pp_1_10 = i_multiplier[1] & i_multiplicand[10];
wire w_pp_1_11 = i_multiplier[1] & i_multiplicand[11];
wire w_pp_1_12 = i_multiplier[1] & i_multiplicand[12];
wire w_pp_1_13 = i_multiplier[1] & i_multiplicand[13];
wire w_pp_1_14 = i_multiplier[1] & i_multiplicand[14];
wire w_pp_1_15 = i_multiplier[1] & i_multiplicand[15];
wire w_pp_2_0 = i_multiplier[2] & i_multiplicand[0];
wire w_pp_2_1 = i_multiplier[2] & i_multiplicand[1];
wire w_pp_2_2 = i_multiplier[2] & i_multiplicand[2];
wire w_pp_2_3 = i_multiplier[2] & i_multiplicand[3];
wire w_pp_2_4 = i_multiplier[2] & i_multiplicand[4];
wire w_pp_2_5 = i_multiplier[2] & i_multiplicand[5];
wire w_pp_2_6 = i_multiplier[2] & i_multiplicand[6];
wire w_pp_2_7 = i_multiplier[2] & i_multiplicand[7];
wire w_pp_2_8 = i_multiplier[2] & i_multiplicand[8];
wire w_pp_2_9 = i_multiplier[2] & i_multiplicand[9];
wire w_pp_2_10 = i_multiplier[2] & i_multiplicand[10];
wire w_pp_2_11 = i_multiplier[2] & i_multiplicand[11];
wire w_pp_2_12 = i_multiplier[2] & i_multiplicand[12];
wire w_pp_2_13 = i_multiplier[2] & i_multiplicand[13];
wire w_pp_2_14 = i_multiplier[2] & i_multiplicand[14];
wire w_pp_2_15 = i_multiplier[2] & i_multiplicand[15];
wire w_pp_3_0 = i_multiplier[3] & i_multiplicand[0];
wire w_pp_3_1 = i_multiplier[3] & i_multiplicand[1];
wire w_pp_3_2 = i_multiplier[3] & i_multiplicand[2];
wire w_pp_3_3 = i_multiplier[3] & i_multiplicand[3];
wire w_pp_3_4 = i_multiplier[3] & i_multiplicand[4];
wire w_pp_3_5 = i_multiplier[3] & i_multiplicand[5];
wire w_pp_3_6 = i_multiplier[3] & i_multiplicand[6];
wire w_pp_3_7 = i_multiplier[3] & i_multiplicand[7];
wire w_pp_3_8 = i_multiplier[3] & i_multiplicand[8];
wire w_pp_3_9 = i_multiplier[3] & i_multiplicand[9];
wire w_pp_3_10 = i_multiplier[3] & i_multiplicand[10];
wire w_pp_3_11 = i_multiplier[3] & i_multiplicand[11];
wire w_pp_3_12 = i_multiplier[3] & i_multiplicand[12];
wire w_pp_3_13 = i_multiplier[3] & i_multiplicand[13];
wire w_pp_3_14 = i_multiplier[3] & i_multiplicand[14];
wire w_pp_3_15 = i_multiplier[3] & i_multiplicand[15];
wire w_pp_4_0 = i_multiplier[4] & i_multiplicand[0];
wire w_pp_4_1 = i_multiplier[4] & i_multiplicand[1];
wire w_pp_4_2 = i_multiplier[4] & i_multiplicand[2];
wire w_pp_4_3 = i_multiplier[4] & i_multiplicand[3];
wire w_pp_4_4 = i_multiplier[4] & i_multiplicand[4];
wire w_pp_4_5 = i_multiplier[4] & i_multiplicand[5];
wire w_pp_4_6 = i_multiplier[4] & i_multiplicand[6];
wire w_pp_4_7 = i_multiplier[4] & i_multiplicand[7];
wire w_pp_4_8 = i_multiplier[4] & i_multiplicand[8];
wire w_pp_4_9 = i_multiplier[4] & i_multiplicand[9];
wire w_pp_4_10 = i_multiplier[4] & i_multiplicand[10];
wire w_pp_4_11 = i_multiplier[4] & i_multiplicand[11];
wire w_pp_4_12 = i_multiplier[4] & i_multiplicand[12];
wire w_pp_4_13 = i_multiplier[4] & i_multiplicand[13];
wire w_pp_4_14 = i_multiplier[4] & i_multiplicand[14];
wire w_pp_4_15 = i_multiplier[4] & i_multiplicand[15];
wire w_pp_5_0 = i_multiplier[5] & i_multiplicand[0];
wire w_pp_5_1 = i_multiplier[5] & i_multiplicand[1];
wire w_pp_5_2 = i_multiplier[5] & i_multiplicand[2];
wire w_pp_5_3 = i_multiplier[5] & i_multiplicand[3];
wire w_pp_5_4 = i_multiplier[5] & i_multiplicand[4];
wire w_pp_5_5 = i_multiplier[5] & i_multiplicand[5];
wire w_pp_5_6 = i_multiplier[5] & i_multiplicand[6];
wire w_pp_5_7 = i_multiplier[5] & i_multiplicand[7];
wire w_pp_5_8 = i_multiplier[5] & i_multiplicand[8];
wire w_pp_5_9 = i_multiplier[5] & i_multiplicand[9];
wire w_pp_5_10 = i_multiplier[5] & i_multiplicand[10];
wire w_pp_5_11 = i_multiplier[5] & i_multiplicand[11];
wire w_pp_5_12 = i_multiplier[5] & i_multiplicand[12];
wire w_pp_5_13 = i_multiplier[5] & i_multiplicand[13];
wire w_pp_5_14 = i_multiplier[5] & i_multiplicand[14];
wire w_pp_5_15 = i_multiplier[5] & i_multiplicand[15];
wire w_pp_6_0 = i_multiplier[6] & i_multiplicand[0];
wire w_pp_6_1 = i_multiplier[6] & i_multiplicand[1];
wire w_pp_6_2 = i_multiplier[6] & i_multiplicand[2];
wire w_pp_6_3 = i_multiplier[6] & i_multiplicand[3];
wire w_pp_6_4 = i_multiplier[6] & i_multiplicand[4];
wire w_pp_6_5 = i_multiplier[6] & i_multiplicand[5];
wire w_pp_6_6 = i_multiplier[6] & i_multiplicand[6];
wire w_pp_6_7 = i_multiplier[6] & i_multiplicand[7];
wire w_pp_6_8 = i_multiplier[6] & i_multiplicand[8];
wire w_pp_6_9 = i_multiplier[6] & i_multiplicand[9];
wire w_pp_6_10 = i_multiplier[6] & i_multiplicand[10];
wire w_pp_6_11 = i_multiplier[6] & i_multiplicand[11];
wire w_pp_6_12 = i_multiplier[6] & i_multiplicand[12];
wire w_pp_6_13 = i_multiplier[6] & i_multiplicand[13];
wire w_pp_6_14 = i_multiplier[6] & i_multiplicand[14];
wire w_pp_6_15 = i_multiplier[6] & i_multiplicand[15];
wire w_pp_7_0 = i_multiplier[7] & i_multiplicand[0];
wire w_pp_7_1 = i_multiplier[7] & i_multiplicand[1];
wire w_pp_7_2 = i_multiplier[7] & i_multiplicand[2];
wire w_pp_7_3 = i_multiplier[7] & i_multiplicand[3];
wire w_pp_7_4 = i_multiplier[7] & i_multiplicand[4];
wire w_pp_7_5 = i_multiplier[7] & i_multiplicand[5];
wire w_pp_7_6 = i_multiplier[7] & i_multiplicand[6];
wire w_pp_7_7 = i_multiplier[7] & i_multiplicand[7];
wire w_pp_7_8 = i_multiplier[7] & i_multiplicand[8];
wire w_pp_7_9 = i_multiplier[7] & i_multiplicand[9];
wire w_pp_7_10 = i_multiplier[7] & i_multiplicand[10];
wire w_pp_7_11 = i_multiplier[7] & i_multiplicand[11];
wire w_pp_7_12 = i_multiplier[7] & i_multiplicand[12];
wire w_pp_7_13 = i_multiplier[7] & i_multiplicand[13];
wire w_pp_7_14 = i_multiplier[7] & i_multiplicand[14];
wire w_pp_7_15 = i_multiplier[7] & i_multiplicand[15];
wire w_pp_8_0 = i_multiplier[8] & i_multiplicand[0];
wire w_pp_8_1 = i_multiplier[8] & i_multiplicand[1];
wire w_pp_8_2 = i_multiplier[8] & i_multiplicand[2];
wire w_pp_8_3 = i_multiplier[8] & i_multiplicand[3];
wire w_pp_8_4 = i_multiplier[8] & i_multiplicand[4];
wire w_pp_8_5 = i_multiplier[8] & i_multiplicand[5];
wire w_pp_8_6 = i_multiplier[8] & i_multiplicand[6];
wire w_pp_8_7 = i_multiplier[8] & i_multiplicand[7];
wire w_pp_8_8 = i_multiplier[8] & i_multiplicand[8];
wire w_pp_8_9 = i_multiplier[8] & i_multiplicand[9];
wire w_pp_8_10 = i_multiplier[8] & i_multiplicand[10];
wire w_pp_8_11 = i_multiplier[8] & i_multiplicand[11];
wire w_pp_8_12 = i_multiplier[8] & i_multiplicand[12];
wire w_pp_8_13 = i_multiplier[8] & i_multiplicand[13];
wire w_pp_8_14 = i_multiplier[8] & i_multiplicand[14];
wire w_pp_8_15 = i_multiplier[8] & i_multiplicand[15];
wire w_pp_9_0 = i_multiplier[9] & i_multiplicand[0];
wire w_pp_9_1 = i_multiplier[9] & i_multiplicand[1];
wire w_pp_9_2 = i_multiplier[9] & i_multiplicand[2];
wire w_pp_9_3 = i_multiplier[9] & i_multiplicand[3];
wire w_pp_9_4 = i_multiplier[9] & i_multiplicand[4];
wire w_pp_9_5 = i_multiplier[9] & i_multiplicand[5];
wire w_pp_9_6 = i_multiplier[9] & i_multiplicand[6];
wire w_pp_9_7 = i_multiplier[9] & i_multiplicand[7];
wire w_pp_9_8 = i_multiplier[9] & i_multiplicand[8];
wire w_pp_9_9 = i_multiplier[9] & i_multiplicand[9];
wire w_pp_9_10 = i_multiplier[9] & i_multiplicand[10];
wire w_pp_9_11 = i_multiplier[9] & i_multiplicand[11];
wire w_pp_9_12 = i_multiplier[9] & i_multiplicand[12];
wire w_pp_9_13 = i_multiplier[9] & i_multiplicand[13];
wire w_pp_9_14 = i_multiplier[9] & i_multiplicand[14];
wire w_pp_9_15 = i_multiplier[9] & i_multiplicand[15];
wire w_pp_10_0 = i_multiplier[10] & i_multiplicand[0];
wire w_pp_10_1 = i_multiplier[10] & i_multiplicand[1];
wire w_pp_10_2 = i_multiplier[10] & i_multiplicand[2];
wire w_pp_10_3 = i_multiplier[10] & i_multiplicand[3];
wire w_pp_10_4 = i_multiplier[10] & i_multiplicand[4];
wire w_pp_10_5 = i_multiplier[10] & i_multiplicand[5];
wire w_pp_10_6 = i_multiplier[10] & i_multiplicand[6];
wire w_pp_10_7 = i_multiplier[10] & i_multiplicand[7];
wire w_pp_10_8 = i_multiplier[10] & i_multiplicand[8];
wire w_pp_10_9 = i_multiplier[10] & i_multiplicand[9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_11_0 = i_multiplier[11] & i_multiplicand[0];
wire w_pp_11_1 = i_multiplier[11] & i_multiplicand[1];
wire w_pp_11_2 = i_multiplier[11] & i_multiplicand[2];
wire w_pp_11_3 = i_multiplier[11] & i_multiplicand[3];
wire w_pp_11_4 = i_multiplier[11] & i_multiplicand[4];
wire w_pp_11_5 = i_multiplier[11] & i_multiplicand[5];
wire w_pp_11_6 = i_multiplier[11] & i_multiplicand[6];
wire w_pp_11_7 = i_multiplier[11] & i_multiplicand[7];
wire w_pp_11_8 = i_multiplier[11] & i_multiplicand[8];
wire w_pp_11_9 = i_multiplier[11] & i_multiplicand[9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_12_0 = i_multiplier[12] & i_multiplicand[0];
wire w_pp_12_1 = i_multiplier[12] & i_multiplicand[1];
wire w_pp_12_2 = i_multiplier[12] & i_multiplicand[2];
wire w_pp_12_3 = i_multiplier[12] & i_multiplicand[3];
wire w_pp_12_4 = i_multiplier[12] & i_multiplicand[4];
wire w_pp_12_5 = i_multiplier[12] & i_multiplicand[5];
wire w_pp_12_6 = i_multiplier[12] & i_multiplicand[6];
wire w_pp_12_7 = i_multiplier[12] & i_multiplicand[7];
wire w_pp_12_8 = i_multiplier[12] & i_multiplicand[8];
wire w_pp_12_9 = i_multiplier[12] & i_multiplicand[9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_13_0 = i_multiplier[13] & i_multiplicand[0];
wire w_pp_13_1 = i_multiplier[13] & i_multiplicand[1];
wire w_pp_13_2 = i_multiplier[13] & i_multiplicand[2];
wire w_pp_13_3 = i_multiplier[13] & i_multiplicand[3];
wire w_pp_13_4 = i_multiplier[13] & i_multiplicand[4];
wire w_pp_13_5 = i_multiplier[13] & i_multiplicand[5];
wire w_pp_13_6 = i_multiplier[13] & i_multiplicand[6];
wire w_pp_13_7 = i_multiplier[13] & i_multiplicand[7];
wire w_pp_13_8 = i_multiplier[13] & i_multiplicand[8];
wire w_pp_13_9 = i_multiplier[13] & i_multiplicand[9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_14_0 = i_multiplier[14] & i_multiplicand[0];
wire w_pp_14_1 = i_multiplier[14] & i_multiplicand[1];
wire w_pp_14_2 = i_multiplier[14] & i_multiplicand[2];
wire w_pp_14_3 = i_multiplier[14] & i_multiplicand[3];
wire w_pp_14_4 = i_multiplier[14] & i_multiplicand[4];
wire w_pp_14_5 = i_multiplier[14] & i_multiplicand[5];
wire w_pp_14_6 = i_multiplier[14] & i_multiplicand[6];
wire w_pp_14_7 = i_multiplier[14] & i_multiplicand[7];
wire w_pp_14_8 = i_multiplier[14] & i_multiplicand[8];
wire w_pp_14_9 = i_multiplier[14] & i_multiplicand[9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_15_0 = i_multiplier[15] & i_multiplicand[0];
wire w_pp_15_1 = i_multiplier[15] & i_multiplicand[1];
wire w_pp_15_2 = i_multiplier[15] & i_multiplicand[2];
wire w_pp_15_3 = i_multiplier[15] & i_multiplicand[3];
wire w_pp_15_4 = i_multiplier[15] & i_multiplicand[4];
wire w_pp_15_5 = i_multiplier[15] & i_multiplicand[5];
wire w_pp_15_6 = i_multiplier[15] & i_multiplicand[6];
wire w_pp_15_7 = i_multiplier[15] & i_multiplicand[7];
wire w_pp_15_8 = i_multiplier[15] & i_multiplicand[8];
wire w_pp_15_9 = i_multiplier[15] & i_multiplicand[9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];

// Partial products reduction using Wallace tree
wire w_sum_1_2, w_carry_1_2;
math_adder_half HA_1_2(.i_a(w_pp_0_1), .i_b(w_pp_1_0), .ow_sum(w_sum_1_2), .ow_c(w_carry_1_2));
wire w_sum_2_4, w_carry_2_4;
math_adder_carry_save CSA_2_4(.i_a(w_pp_0_2), .i_b(w_pp_1_1), .i_c(w_pp_2_0), .ow_sum(w_sum_2_4), .ow_c(w_carry_2_4));
wire w_sum_2_2, w_carry_2_2;
math_adder_half HA_2_2(.i_a(w_carry_1_2), .i_b(w_sum_2_4), .ow_sum(w_sum_2_2), .ow_c(w_carry_2_2));
wire w_sum_3_6, w_carry_3_6;
math_adder_carry_save CSA_3_6(.i_a(w_pp_0_3), .i_b(w_pp_1_2), .i_c(w_pp_2_1), .ow_sum(w_sum_3_6), .ow_c(w_carry_3_6));
wire w_sum_3_4, w_carry_3_4;
math_adder_carry_save CSA_3_4(.i_a(w_pp_3_0), .i_b(w_carry_2_4), .i_c(w_carry_2_2), .ow_sum(w_sum_3_4), .ow_c(w_carry_3_4));
wire w_sum_3_2, w_carry_3_2;
math_adder_half HA_3_2(.i_a(w_sum_3_6), .i_b(w_sum_3_4), .ow_sum(w_sum_3_2), .ow_c(w_carry_3_2));
wire w_sum_4_8, w_carry_4_8;
math_adder_carry_save CSA_4_8(.i_a(w_pp_0_4), .i_b(w_pp_1_3), .i_c(w_pp_2_2), .ow_sum(w_sum_4_8), .ow_c(w_carry_4_8));
wire w_sum_4_6, w_carry_4_6;
math_adder_carry_save CSA_4_6(.i_a(w_pp_3_1), .i_b(w_pp_4_0), .i_c(w_carry_3_6), .ow_sum(w_sum_4_6), .ow_c(w_carry_4_6));
wire w_sum_4_4, w_carry_4_4;
math_adder_carry_save CSA_4_4(.i_a(w_carry_3_4), .i_b(w_carry_3_2), .i_c(w_sum_4_8), .ow_sum(w_sum_4_4), .ow_c(w_carry_4_4));
wire w_sum_4_2, w_carry_4_2;
math_adder_half HA_4_2(.i_a(w_sum_4_6), .i_b(w_sum_4_4), .ow_sum(w_sum_4_2), .ow_c(w_carry_4_2));
wire w_sum_5_10, w_carry_5_10;
math_adder_carry_save CSA_5_10(.i_a(w_pp_0_5), .i_b(w_pp_1_4), .i_c(w_pp_2_3), .ow_sum(w_sum_5_10), .ow_c(w_carry_5_10));
wire w_sum_5_8, w_carry_5_8;
math_adder_carry_save CSA_5_8(.i_a(w_pp_3_2), .i_b(w_pp_4_1), .i_c(w_pp_5_0), .ow_sum(w_sum_5_8), .ow_c(w_carry_5_8));
wire w_sum_5_6, w_carry_5_6;
math_adder_carry_save CSA_5_6(.i_a(w_carry_4_8), .i_b(w_carry_4_6), .i_c(w_carry_4_4), .ow_sum(w_sum_5_6), .ow_c(w_carry_5_6));
wire w_sum_5_4, w_carry_5_4;
math_adder_carry_save CSA_5_4(.i_a(w_carry_4_2), .i_b(w_sum_5_10), .i_c(w_sum_5_8), .ow_sum(w_sum_5_4), .ow_c(w_carry_5_4));
wire w_sum_5_2, w_carry_5_2;
math_adder_half HA_5_2(.i_a(w_sum_5_6), .i_b(w_sum_5_4), .ow_sum(w_sum_5_2), .ow_c(w_carry_5_2));
wire w_sum_6_12, w_carry_6_12;
math_adder_carry_save CSA_6_12(.i_a(w_pp_0_6), .i_b(w_pp_1_5), .i_c(w_pp_2_4), .ow_sum(w_sum_6_12), .ow_c(w_carry_6_12));
wire w_sum_6_10, w_carry_6_10;
math_adder_carry_save CSA_6_10(.i_a(w_pp_3_3), .i_b(w_pp_4_2), .i_c(w_pp_5_1), .ow_sum(w_sum_6_10), .ow_c(w_carry_6_10));
wire w_sum_6_8, w_carry_6_8;
math_adder_carry_save CSA_6_8(.i_a(w_pp_6_0), .i_b(w_carry_5_10), .i_c(w_carry_5_8), .ow_sum(w_sum_6_8), .ow_c(w_carry_6_8));
wire w_sum_6_6, w_carry_6_6;
math_adder_carry_save CSA_6_6(.i_a(w_carry_5_6), .i_b(w_carry_5_4), .i_c(w_carry_5_2), .ow_sum(w_sum_6_6), .ow_c(w_carry_6_6));
wire w_sum_6_4, w_carry_6_4;
math_adder_carry_save CSA_6_4(.i_a(w_sum_6_12), .i_b(w_sum_6_10), .i_c(w_sum_6_8), .ow_sum(w_sum_6_4), .ow_c(w_carry_6_4));
wire w_sum_6_2, w_carry_6_2;
math_adder_half HA_6_2(.i_a(w_sum_6_6), .i_b(w_sum_6_4), .ow_sum(w_sum_6_2), .ow_c(w_carry_6_2));
wire w_sum_7_14, w_carry_7_14;
math_adder_carry_save CSA_7_14(.i_a(w_pp_0_7), .i_b(w_pp_1_6), .i_c(w_pp_2_5), .ow_sum(w_sum_7_14), .ow_c(w_carry_7_14));
wire w_sum_7_12, w_carry_7_12;
math_adder_carry_save CSA_7_12(.i_a(w_pp_3_4), .i_b(w_pp_4_3), .i_c(w_pp_5_2), .ow_sum(w_sum_7_12), .ow_c(w_carry_7_12));
wire w_sum_7_10, w_carry_7_10;
math_adder_carry_save CSA_7_10(.i_a(w_pp_6_1), .i_b(w_pp_7_0), .i_c(w_carry_6_12), .ow_sum(w_sum_7_10), .ow_c(w_carry_7_10));
wire w_sum_7_8, w_carry_7_8;
math_adder_carry_save CSA_7_8(.i_a(w_carry_6_10), .i_b(w_carry_6_8), .i_c(w_carry_6_6), .ow_sum(w_sum_7_8), .ow_c(w_carry_7_8));
wire w_sum_7_6, w_carry_7_6;
math_adder_carry_save CSA_7_6(.i_a(w_carry_6_4), .i_b(w_carry_6_2), .i_c(w_sum_7_14), .ow_sum(w_sum_7_6), .ow_c(w_carry_7_6));
wire w_sum_7_4, w_carry_7_4;
math_adder_carry_save CSA_7_4(.i_a(w_sum_7_12), .i_b(w_sum_7_10), .i_c(w_sum_7_8), .ow_sum(w_sum_7_4), .ow_c(w_carry_7_4));
wire w_sum_7_2, w_carry_7_2;
math_adder_half HA_7_2(.i_a(w_sum_7_6), .i_b(w_sum_7_4), .ow_sum(w_sum_7_2), .ow_c(w_carry_7_2));
wire w_sum_8_16, w_carry_8_16;
math_adder_carry_save CSA_8_16(.i_a(w_pp_0_8), .i_b(w_pp_1_7), .i_c(w_pp_2_6), .ow_sum(w_sum_8_16), .ow_c(w_carry_8_16));
wire w_sum_8_14, w_carry_8_14;
math_adder_carry_save CSA_8_14(.i_a(w_pp_3_5), .i_b(w_pp_4_4), .i_c(w_pp_5_3), .ow_sum(w_sum_8_14), .ow_c(w_carry_8_14));
wire w_sum_8_12, w_carry_8_12;
math_adder_carry_save CSA_8_12(.i_a(w_pp_6_2), .i_b(w_pp_7_1), .i_c(w_pp_8_0), .ow_sum(w_sum_8_12), .ow_c(w_carry_8_12));
wire w_sum_8_10, w_carry_8_10;
math_adder_carry_save CSA_8_10(.i_a(w_carry_7_14), .i_b(w_carry_7_12), .i_c(w_carry_7_10), .ow_sum(w_sum_8_10), .ow_c(w_carry_8_10));
wire w_sum_8_8, w_carry_8_8;
math_adder_carry_save CSA_8_8(.i_a(w_carry_7_8), .i_b(w_carry_7_6), .i_c(w_carry_7_4), .ow_sum(w_sum_8_8), .ow_c(w_carry_8_8));
wire w_sum_8_6, w_carry_8_6;
math_adder_carry_save CSA_8_6(.i_a(w_carry_7_2), .i_b(w_sum_8_16), .i_c(w_sum_8_14), .ow_sum(w_sum_8_6), .ow_c(w_carry_8_6));
wire w_sum_8_4, w_carry_8_4;
math_adder_carry_save CSA_8_4(.i_a(w_sum_8_12), .i_b(w_sum_8_10), .i_c(w_sum_8_8), .ow_sum(w_sum_8_4), .ow_c(w_carry_8_4));
wire w_sum_8_2, w_carry_8_2;
math_adder_half HA_8_2(.i_a(w_sum_8_6), .i_b(w_sum_8_4), .ow_sum(w_sum_8_2), .ow_c(w_carry_8_2));
wire w_sum_9_18, w_carry_9_18;
math_adder_carry_save CSA_9_18(.i_a(w_pp_0_9), .i_b(w_pp_1_8), .i_c(w_pp_2_7), .ow_sum(w_sum_9_18), .ow_c(w_carry_9_18));
wire w_sum_9_16, w_carry_9_16;
math_adder_carry_save CSA_9_16(.i_a(w_pp_3_6), .i_b(w_pp_4_5), .i_c(w_pp_5_4), .ow_sum(w_sum_9_16), .ow_c(w_carry_9_16));
wire w_sum_9_14, w_carry_9_14;
math_adder_carry_save CSA_9_14(.i_a(w_pp_6_3), .i_b(w_pp_7_2), .i_c(w_pp_8_1), .ow_sum(w_sum_9_14), .ow_c(w_carry_9_14));
wire w_sum_9_12, w_carry_9_12;
math_adder_carry_save CSA_9_12(.i_a(w_pp_9_0), .i_b(w_carry_8_16), .i_c(w_carry_8_14), .ow_sum(w_sum_9_12), .ow_c(w_carry_9_12));
wire w_sum_9_10, w_carry_9_10;
math_adder_carry_save CSA_9_10(.i_a(w_carry_8_12), .i_b(w_carry_8_10), .i_c(w_carry_8_8), .ow_sum(w_sum_9_10), .ow_c(w_carry_9_10));
wire w_sum_9_8, w_carry_9_8;
math_adder_carry_save CSA_9_8(.i_a(w_carry_8_6), .i_b(w_carry_8_4), .i_c(w_carry_8_2), .ow_sum(w_sum_9_8), .ow_c(w_carry_9_8));
wire w_sum_9_6, w_carry_9_6;
math_adder_carry_save CSA_9_6(.i_a(w_sum_9_18), .i_b(w_sum_9_16), .i_c(w_sum_9_14), .ow_sum(w_sum_9_6), .ow_c(w_carry_9_6));
wire w_sum_9_4, w_carry_9_4;
math_adder_carry_save CSA_9_4(.i_a(w_sum_9_12), .i_b(w_sum_9_10), .i_c(w_sum_9_8), .ow_sum(w_sum_9_4), .ow_c(w_carry_9_4));
wire w_sum_9_2, w_carry_9_2;
math_adder_half HA_9_2(.i_a(w_sum_9_6), .i_b(w_sum_9_4), .ow_sum(w_sum_9_2), .ow_c(w_carry_9_2));
wire w_sum_10_20, w_carry_10_20;
math_adder_carry_save CSA_10_20(.i_a(w_pp_0_10), .i_b(w_pp_1_9), .i_c(w_pp_2_8), .ow_sum(w_sum_10_20), .ow_c(w_carry_10_20));
wire w_sum_10_18, w_carry_10_18;
math_adder_carry_save CSA_10_18(.i_a(w_pp_3_7), .i_b(w_pp_4_6), .i_c(w_pp_5_5), .ow_sum(w_sum_10_18), .ow_c(w_carry_10_18));
wire w_sum_10_16, w_carry_10_16;
math_adder_carry_save CSA_10_16(.i_a(w_pp_6_4), .i_b(w_pp_7_3), .i_c(w_pp_8_2), .ow_sum(w_sum_10_16), .ow_c(w_carry_10_16));
wire w_sum_10_14, w_carry_10_14;
math_adder_carry_save CSA_10_14(.i_a(w_pp_9_1), .i_b(w_pp_10_0), .i_c(w_carry_9_18), .ow_sum(w_sum_10_14), .ow_c(w_carry_10_14));
wire w_sum_10_12, w_carry_10_12;
math_adder_carry_save CSA_10_12(.i_a(w_carry_9_16), .i_b(w_carry_9_14), .i_c(w_carry_9_12), .ow_sum(w_sum_10_12), .ow_c(w_carry_10_12));
wire w_sum_10_10, w_carry_10_10;
math_adder_carry_save CSA_10_10(.i_a(w_carry_9_10), .i_b(w_carry_9_8), .i_c(w_carry_9_6), .ow_sum(w_sum_10_10), .ow_c(w_carry_10_10));
wire w_sum_10_8, w_carry_10_8;
math_adder_carry_save CSA_10_8(.i_a(w_carry_9_4), .i_b(w_carry_9_2), .i_c(w_sum_10_20), .ow_sum(w_sum_10_8), .ow_c(w_carry_10_8));
wire w_sum_10_6, w_carry_10_6;
math_adder_carry_save CSA_10_6(.i_a(w_sum_10_18), .i_b(w_sum_10_16), .i_c(w_sum_10_14), .ow_sum(w_sum_10_6), .ow_c(w_carry_10_6));
wire w_sum_10_4, w_carry_10_4;
math_adder_carry_save CSA_10_4(.i_a(w_sum_10_12), .i_b(w_sum_10_10), .i_c(w_sum_10_8), .ow_sum(w_sum_10_4), .ow_c(w_carry_10_4));
wire w_sum_10_2, w_carry_10_2;
math_adder_half HA_10_2(.i_a(w_sum_10_6), .i_b(w_sum_10_4), .ow_sum(w_sum_10_2), .ow_c(w_carry_10_2));
wire w_sum_11_22, w_carry_11_22;
math_adder_carry_save CSA_11_22(.i_a(w_pp_0_11), .i_b(w_pp_1_10), .i_c(w_pp_2_9), .ow_sum(w_sum_11_22), .ow_c(w_carry_11_22));
wire w_sum_11_20, w_carry_11_20;
math_adder_carry_save CSA_11_20(.i_a(w_pp_3_8), .i_b(w_pp_4_7), .i_c(w_pp_5_6), .ow_sum(w_sum_11_20), .ow_c(w_carry_11_20));
wire w_sum_11_18, w_carry_11_18;
math_adder_carry_save CSA_11_18(.i_a(w_pp_6_5), .i_b(w_pp_7_4), .i_c(w_pp_8_3), .ow_sum(w_sum_11_18), .ow_c(w_carry_11_18));
wire w_sum_11_16, w_carry_11_16;
math_adder_carry_save CSA_11_16(.i_a(w_pp_9_2), .i_b(w_pp_10_1), .i_c(w_pp_11_0), .ow_sum(w_sum_11_16), .ow_c(w_carry_11_16));
wire w_sum_11_14, w_carry_11_14;
math_adder_carry_save CSA_11_14(.i_a(w_carry_10_20), .i_b(w_carry_10_18), .i_c(w_carry_10_16), .ow_sum(w_sum_11_14), .ow_c(w_carry_11_14));
wire w_sum_11_12, w_carry_11_12;
math_adder_carry_save CSA_11_12(.i_a(w_carry_10_14), .i_b(w_carry_10_12), .i_c(w_carry_10_10), .ow_sum(w_sum_11_12), .ow_c(w_carry_11_12));
wire w_sum_11_10, w_carry_11_10;
math_adder_carry_save CSA_11_10(.i_a(w_carry_10_8), .i_b(w_carry_10_6), .i_c(w_carry_10_4), .ow_sum(w_sum_11_10), .ow_c(w_carry_11_10));
wire w_sum_11_8, w_carry_11_8;
math_adder_carry_save CSA_11_8(.i_a(w_carry_10_2), .i_b(w_sum_11_22), .i_c(w_sum_11_20), .ow_sum(w_sum_11_8), .ow_c(w_carry_11_8));
wire w_sum_11_6, w_carry_11_6;
math_adder_carry_save CSA_11_6(.i_a(w_sum_11_18), .i_b(w_sum_11_16), .i_c(w_sum_11_14), .ow_sum(w_sum_11_6), .ow_c(w_carry_11_6));
wire w_sum_11_4, w_carry_11_4;
math_adder_carry_save CSA_11_4(.i_a(w_sum_11_12), .i_b(w_sum_11_10), .i_c(w_sum_11_8), .ow_sum(w_sum_11_4), .ow_c(w_carry_11_4));
wire w_sum_11_2, w_carry_11_2;
math_adder_half HA_11_2(.i_a(w_sum_11_6), .i_b(w_sum_11_4), .ow_sum(w_sum_11_2), .ow_c(w_carry_11_2));
wire w_sum_12_24, w_carry_12_24;
math_adder_carry_save CSA_12_24(.i_a(w_pp_0_12), .i_b(w_pp_1_11), .i_c(w_pp_2_10), .ow_sum(w_sum_12_24), .ow_c(w_carry_12_24));
wire w_sum_12_22, w_carry_12_22;
math_adder_carry_save CSA_12_22(.i_a(w_pp_3_9), .i_b(w_pp_4_8), .i_c(w_pp_5_7), .ow_sum(w_sum_12_22), .ow_c(w_carry_12_22));
wire w_sum_12_20, w_carry_12_20;
math_adder_carry_save CSA_12_20(.i_a(w_pp_6_6), .i_b(w_pp_7_5), .i_c(w_pp_8_4), .ow_sum(w_sum_12_20), .ow_c(w_carry_12_20));
wire w_sum_12_18, w_carry_12_18;
math_adder_carry_save CSA_12_18(.i_a(w_pp_9_3), .i_b(w_pp_10_2), .i_c(w_pp_11_1), .ow_sum(w_sum_12_18), .ow_c(w_carry_12_18));
wire w_sum_12_16, w_carry_12_16;
math_adder_carry_save CSA_12_16(.i_a(w_pp_12_0), .i_b(w_carry_11_22), .i_c(w_carry_11_20), .ow_sum(w_sum_12_16), .ow_c(w_carry_12_16));
wire w_sum_12_14, w_carry_12_14;
math_adder_carry_save CSA_12_14(.i_a(w_carry_11_18), .i_b(w_carry_11_16), .i_c(w_carry_11_14), .ow_sum(w_sum_12_14), .ow_c(w_carry_12_14));
wire w_sum_12_12, w_carry_12_12;
math_adder_carry_save CSA_12_12(.i_a(w_carry_11_12), .i_b(w_carry_11_10), .i_c(w_carry_11_8), .ow_sum(w_sum_12_12), .ow_c(w_carry_12_12));
wire w_sum_12_10, w_carry_12_10;
math_adder_carry_save CSA_12_10(.i_a(w_carry_11_6), .i_b(w_carry_11_4), .i_c(w_carry_11_2), .ow_sum(w_sum_12_10), .ow_c(w_carry_12_10));
wire w_sum_12_8, w_carry_12_8;
math_adder_carry_save CSA_12_8(.i_a(w_sum_12_24), .i_b(w_sum_12_22), .i_c(w_sum_12_20), .ow_sum(w_sum_12_8), .ow_c(w_carry_12_8));
wire w_sum_12_6, w_carry_12_6;
math_adder_carry_save CSA_12_6(.i_a(w_sum_12_18), .i_b(w_sum_12_16), .i_c(w_sum_12_14), .ow_sum(w_sum_12_6), .ow_c(w_carry_12_6));
wire w_sum_12_4, w_carry_12_4;
math_adder_carry_save CSA_12_4(.i_a(w_sum_12_12), .i_b(w_sum_12_10), .i_c(w_sum_12_8), .ow_sum(w_sum_12_4), .ow_c(w_carry_12_4));
wire w_sum_12_2, w_carry_12_2;
math_adder_half HA_12_2(.i_a(w_sum_12_6), .i_b(w_sum_12_4), .ow_sum(w_sum_12_2), .ow_c(w_carry_12_2));
wire w_sum_13_26, w_carry_13_26;
math_adder_carry_save CSA_13_26(.i_a(w_pp_0_13), .i_b(w_pp_1_12), .i_c(w_pp_2_11), .ow_sum(w_sum_13_26), .ow_c(w_carry_13_26));
wire w_sum_13_24, w_carry_13_24;
math_adder_carry_save CSA_13_24(.i_a(w_pp_3_10), .i_b(w_pp_4_9), .i_c(w_pp_5_8), .ow_sum(w_sum_13_24), .ow_c(w_carry_13_24));
wire w_sum_13_22, w_carry_13_22;
math_adder_carry_save CSA_13_22(.i_a(w_pp_6_7), .i_b(w_pp_7_6), .i_c(w_pp_8_5), .ow_sum(w_sum_13_22), .ow_c(w_carry_13_22));
wire w_sum_13_20, w_carry_13_20;
math_adder_carry_save CSA_13_20(.i_a(w_pp_9_4), .i_b(w_pp_10_3), .i_c(w_pp_11_2), .ow_sum(w_sum_13_20), .ow_c(w_carry_13_20));
wire w_sum_13_18, w_carry_13_18;
math_adder_carry_save CSA_13_18(.i_a(w_pp_12_1), .i_b(w_pp_13_0), .i_c(w_carry_12_24), .ow_sum(w_sum_13_18), .ow_c(w_carry_13_18));
wire w_sum_13_16, w_carry_13_16;
math_adder_carry_save CSA_13_16(.i_a(w_carry_12_22), .i_b(w_carry_12_20), .i_c(w_carry_12_18), .ow_sum(w_sum_13_16), .ow_c(w_carry_13_16));
wire w_sum_13_14, w_carry_13_14;
math_adder_carry_save CSA_13_14(.i_a(w_carry_12_16), .i_b(w_carry_12_14), .i_c(w_carry_12_12), .ow_sum(w_sum_13_14), .ow_c(w_carry_13_14));
wire w_sum_13_12, w_carry_13_12;
math_adder_carry_save CSA_13_12(.i_a(w_carry_12_10), .i_b(w_carry_12_8), .i_c(w_carry_12_6), .ow_sum(w_sum_13_12), .ow_c(w_carry_13_12));
wire w_sum_13_10, w_carry_13_10;
math_adder_carry_save CSA_13_10(.i_a(w_carry_12_4), .i_b(w_carry_12_2), .i_c(w_sum_13_26), .ow_sum(w_sum_13_10), .ow_c(w_carry_13_10));
wire w_sum_13_8, w_carry_13_8;
math_adder_carry_save CSA_13_8(.i_a(w_sum_13_24), .i_b(w_sum_13_22), .i_c(w_sum_13_20), .ow_sum(w_sum_13_8), .ow_c(w_carry_13_8));
wire w_sum_13_6, w_carry_13_6;
math_adder_carry_save CSA_13_6(.i_a(w_sum_13_18), .i_b(w_sum_13_16), .i_c(w_sum_13_14), .ow_sum(w_sum_13_6), .ow_c(w_carry_13_6));
wire w_sum_13_4, w_carry_13_4;
math_adder_carry_save CSA_13_4(.i_a(w_sum_13_12), .i_b(w_sum_13_10), .i_c(w_sum_13_8), .ow_sum(w_sum_13_4), .ow_c(w_carry_13_4));
wire w_sum_13_2, w_carry_13_2;
math_adder_half HA_13_2(.i_a(w_sum_13_6), .i_b(w_sum_13_4), .ow_sum(w_sum_13_2), .ow_c(w_carry_13_2));
wire w_sum_14_28, w_carry_14_28;
math_adder_carry_save CSA_14_28(.i_a(w_pp_0_14), .i_b(w_pp_1_13), .i_c(w_pp_2_12), .ow_sum(w_sum_14_28), .ow_c(w_carry_14_28));
wire w_sum_14_26, w_carry_14_26;
math_adder_carry_save CSA_14_26(.i_a(w_pp_3_11), .i_b(w_pp_4_10), .i_c(w_pp_5_9), .ow_sum(w_sum_14_26), .ow_c(w_carry_14_26));
wire w_sum_14_24, w_carry_14_24;
math_adder_carry_save CSA_14_24(.i_a(w_pp_6_8), .i_b(w_pp_7_7), .i_c(w_pp_8_6), .ow_sum(w_sum_14_24), .ow_c(w_carry_14_24));
wire w_sum_14_22, w_carry_14_22;
math_adder_carry_save CSA_14_22(.i_a(w_pp_9_5), .i_b(w_pp_10_4), .i_c(w_pp_11_3), .ow_sum(w_sum_14_22), .ow_c(w_carry_14_22));
wire w_sum_14_20, w_carry_14_20;
math_adder_carry_save CSA_14_20(.i_a(w_pp_12_2), .i_b(w_pp_13_1), .i_c(w_pp_14_0), .ow_sum(w_sum_14_20), .ow_c(w_carry_14_20));
wire w_sum_14_18, w_carry_14_18;
math_adder_carry_save CSA_14_18(.i_a(w_carry_13_26), .i_b(w_carry_13_24), .i_c(w_carry_13_22), .ow_sum(w_sum_14_18), .ow_c(w_carry_14_18));
wire w_sum_14_16, w_carry_14_16;
math_adder_carry_save CSA_14_16(.i_a(w_carry_13_20), .i_b(w_carry_13_18), .i_c(w_carry_13_16), .ow_sum(w_sum_14_16), .ow_c(w_carry_14_16));
wire w_sum_14_14, w_carry_14_14;
math_adder_carry_save CSA_14_14(.i_a(w_carry_13_14), .i_b(w_carry_13_12), .i_c(w_carry_13_10), .ow_sum(w_sum_14_14), .ow_c(w_carry_14_14));
wire w_sum_14_12, w_carry_14_12;
math_adder_carry_save CSA_14_12(.i_a(w_carry_13_8), .i_b(w_carry_13_6), .i_c(w_carry_13_4), .ow_sum(w_sum_14_12), .ow_c(w_carry_14_12));
wire w_sum_14_10, w_carry_14_10;
math_adder_carry_save CSA_14_10(.i_a(w_carry_13_2), .i_b(w_sum_14_28), .i_c(w_sum_14_26), .ow_sum(w_sum_14_10), .ow_c(w_carry_14_10));
wire w_sum_14_8, w_carry_14_8;
math_adder_carry_save CSA_14_8(.i_a(w_sum_14_24), .i_b(w_sum_14_22), .i_c(w_sum_14_20), .ow_sum(w_sum_14_8), .ow_c(w_carry_14_8));
wire w_sum_14_6, w_carry_14_6;
math_adder_carry_save CSA_14_6(.i_a(w_sum_14_18), .i_b(w_sum_14_16), .i_c(w_sum_14_14), .ow_sum(w_sum_14_6), .ow_c(w_carry_14_6));
wire w_sum_14_4, w_carry_14_4;
math_adder_carry_save CSA_14_4(.i_a(w_sum_14_12), .i_b(w_sum_14_10), .i_c(w_sum_14_8), .ow_sum(w_sum_14_4), .ow_c(w_carry_14_4));
wire w_sum_14_2, w_carry_14_2;
math_adder_half HA_14_2(.i_a(w_sum_14_6), .i_b(w_sum_14_4), .ow_sum(w_sum_14_2), .ow_c(w_carry_14_2));
wire w_sum_15_30, w_carry_15_30;
math_adder_carry_save CSA_15_30(.i_a(w_pp_0_15), .i_b(w_pp_1_14), .i_c(w_pp_2_13), .ow_sum(w_sum_15_30), .ow_c(w_carry_15_30));
wire w_sum_15_28, w_carry_15_28;
math_adder_carry_save CSA_15_28(.i_a(w_pp_3_12), .i_b(w_pp_4_11), .i_c(w_pp_5_10), .ow_sum(w_sum_15_28), .ow_c(w_carry_15_28));
wire w_sum_15_26, w_carry_15_26;
math_adder_carry_save CSA_15_26(.i_a(w_pp_6_9), .i_b(w_pp_7_8), .i_c(w_pp_8_7), .ow_sum(w_sum_15_26), .ow_c(w_carry_15_26));
wire w_sum_15_24, w_carry_15_24;
math_adder_carry_save CSA_15_24(.i_a(w_pp_9_6), .i_b(w_pp_10_5), .i_c(w_pp_11_4), .ow_sum(w_sum_15_24), .ow_c(w_carry_15_24));
wire w_sum_15_22, w_carry_15_22;
math_adder_carry_save CSA_15_22(.i_a(w_pp_12_3), .i_b(w_pp_13_2), .i_c(w_pp_14_1), .ow_sum(w_sum_15_22), .ow_c(w_carry_15_22));
wire w_sum_15_20, w_carry_15_20;
math_adder_carry_save CSA_15_20(.i_a(w_pp_15_0), .i_b(w_carry_14_28), .i_c(w_carry_14_26), .ow_sum(w_sum_15_20), .ow_c(w_carry_15_20));
wire w_sum_15_18, w_carry_15_18;
math_adder_carry_save CSA_15_18(.i_a(w_carry_14_24), .i_b(w_carry_14_22), .i_c(w_carry_14_20), .ow_sum(w_sum_15_18), .ow_c(w_carry_15_18));
wire w_sum_15_16, w_carry_15_16;
math_adder_carry_save CSA_15_16(.i_a(w_carry_14_18), .i_b(w_carry_14_16), .i_c(w_carry_14_14), .ow_sum(w_sum_15_16), .ow_c(w_carry_15_16));
wire w_sum_15_14, w_carry_15_14;
math_adder_carry_save CSA_15_14(.i_a(w_carry_14_12), .i_b(w_carry_14_10), .i_c(w_carry_14_8), .ow_sum(w_sum_15_14), .ow_c(w_carry_15_14));
wire w_sum_15_12, w_carry_15_12;
math_adder_carry_save CSA_15_12(.i_a(w_carry_14_6), .i_b(w_carry_14_4), .i_c(w_carry_14_2), .ow_sum(w_sum_15_12), .ow_c(w_carry_15_12));
wire w_sum_15_10, w_carry_15_10;
math_adder_carry_save CSA_15_10(.i_a(w_sum_15_30), .i_b(w_sum_15_28), .i_c(w_sum_15_26), .ow_sum(w_sum_15_10), .ow_c(w_carry_15_10));
wire w_sum_15_8, w_carry_15_8;
math_adder_carry_save CSA_15_8(.i_a(w_sum_15_24), .i_b(w_sum_15_22), .i_c(w_sum_15_20), .ow_sum(w_sum_15_8), .ow_c(w_carry_15_8));
wire w_sum_15_6, w_carry_15_6;
math_adder_carry_save CSA_15_6(.i_a(w_sum_15_18), .i_b(w_sum_15_16), .i_c(w_sum_15_14), .ow_sum(w_sum_15_6), .ow_c(w_carry_15_6));
wire w_sum_15_4, w_carry_15_4;
math_adder_carry_save CSA_15_4(.i_a(w_sum_15_12), .i_b(w_sum_15_10), .i_c(w_sum_15_8), .ow_sum(w_sum_15_4), .ow_c(w_carry_15_4));
wire w_sum_15_2, w_carry_15_2;
math_adder_half HA_15_2(.i_a(w_sum_15_6), .i_b(w_sum_15_4), .ow_sum(w_sum_15_2), .ow_c(w_carry_15_2));
wire w_sum_16_30, w_carry_16_30;
math_adder_carry_save CSA_16_30(.i_a(w_pp_1_15), .i_b(w_pp_2_14), .i_c(w_pp_3_13), .ow_sum(w_sum_16_30), .ow_c(w_carry_16_30));
wire w_sum_16_28, w_carry_16_28;
math_adder_carry_save CSA_16_28(.i_a(w_pp_4_12), .i_b(w_pp_5_11), .i_c(w_pp_6_10), .ow_sum(w_sum_16_28), .ow_c(w_carry_16_28));
wire w_sum_16_26, w_carry_16_26;
math_adder_carry_save CSA_16_26(.i_a(w_pp_7_9), .i_b(w_pp_8_8), .i_c(w_pp_9_7), .ow_sum(w_sum_16_26), .ow_c(w_carry_16_26));
wire w_sum_16_24, w_carry_16_24;
math_adder_carry_save CSA_16_24(.i_a(w_pp_10_6), .i_b(w_pp_11_5), .i_c(w_pp_12_4), .ow_sum(w_sum_16_24), .ow_c(w_carry_16_24));
wire w_sum_16_22, w_carry_16_22;
math_adder_carry_save CSA_16_22(.i_a(w_pp_13_3), .i_b(w_pp_14_2), .i_c(w_pp_15_1), .ow_sum(w_sum_16_22), .ow_c(w_carry_16_22));
wire w_sum_16_20, w_carry_16_20;
math_adder_carry_save CSA_16_20(.i_a(w_carry_15_30), .i_b(w_carry_15_28), .i_c(w_carry_15_26), .ow_sum(w_sum_16_20), .ow_c(w_carry_16_20));
wire w_sum_16_18, w_carry_16_18;
math_adder_carry_save CSA_16_18(.i_a(w_carry_15_24), .i_b(w_carry_15_22), .i_c(w_carry_15_20), .ow_sum(w_sum_16_18), .ow_c(w_carry_16_18));
wire w_sum_16_16, w_carry_16_16;
math_adder_carry_save CSA_16_16(.i_a(w_carry_15_18), .i_b(w_carry_15_16), .i_c(w_carry_15_14), .ow_sum(w_sum_16_16), .ow_c(w_carry_16_16));
wire w_sum_16_14, w_carry_16_14;
math_adder_carry_save CSA_16_14(.i_a(w_carry_15_12), .i_b(w_carry_15_10), .i_c(w_carry_15_8), .ow_sum(w_sum_16_14), .ow_c(w_carry_16_14));
wire w_sum_16_12, w_carry_16_12;
math_adder_carry_save CSA_16_12(.i_a(w_carry_15_6), .i_b(w_carry_15_4), .i_c(w_carry_15_2), .ow_sum(w_sum_16_12), .ow_c(w_carry_16_12));
wire w_sum_16_10, w_carry_16_10;
math_adder_carry_save CSA_16_10(.i_a(w_sum_16_30), .i_b(w_sum_16_28), .i_c(w_sum_16_26), .ow_sum(w_sum_16_10), .ow_c(w_carry_16_10));
wire w_sum_16_8, w_carry_16_8;
math_adder_carry_save CSA_16_8(.i_a(w_sum_16_24), .i_b(w_sum_16_22), .i_c(w_sum_16_20), .ow_sum(w_sum_16_8), .ow_c(w_carry_16_8));
wire w_sum_16_6, w_carry_16_6;
math_adder_carry_save CSA_16_6(.i_a(w_sum_16_18), .i_b(w_sum_16_16), .i_c(w_sum_16_14), .ow_sum(w_sum_16_6), .ow_c(w_carry_16_6));
wire w_sum_16_4, w_carry_16_4;
math_adder_carry_save CSA_16_4(.i_a(w_sum_16_12), .i_b(w_sum_16_10), .i_c(w_sum_16_8), .ow_sum(w_sum_16_4), .ow_c(w_carry_16_4));
wire w_sum_16_2, w_carry_16_2;
math_adder_half HA_16_2(.i_a(w_sum_16_6), .i_b(w_sum_16_4), .ow_sum(w_sum_16_2), .ow_c(w_carry_16_2));
wire w_sum_17_29, w_carry_17_29;
math_adder_carry_save CSA_17_29(.i_a(w_pp_2_15), .i_b(w_pp_3_14), .i_c(w_pp_4_13), .ow_sum(w_sum_17_29), .ow_c(w_carry_17_29));
wire w_sum_17_27, w_carry_17_27;
math_adder_carry_save CSA_17_27(.i_a(w_pp_5_12), .i_b(w_pp_6_11), .i_c(w_pp_7_10), .ow_sum(w_sum_17_27), .ow_c(w_carry_17_27));
wire w_sum_17_25, w_carry_17_25;
math_adder_carry_save CSA_17_25(.i_a(w_pp_8_9), .i_b(w_pp_9_8), .i_c(w_pp_10_7), .ow_sum(w_sum_17_25), .ow_c(w_carry_17_25));
wire w_sum_17_23, w_carry_17_23;
math_adder_carry_save CSA_17_23(.i_a(w_pp_11_6), .i_b(w_pp_12_5), .i_c(w_pp_13_4), .ow_sum(w_sum_17_23), .ow_c(w_carry_17_23));
wire w_sum_17_21, w_carry_17_21;
math_adder_carry_save CSA_17_21(.i_a(w_pp_14_3), .i_b(w_pp_15_2), .i_c(w_carry_16_30), .ow_sum(w_sum_17_21), .ow_c(w_carry_17_21));
wire w_sum_17_19, w_carry_17_19;
math_adder_carry_save CSA_17_19(.i_a(w_carry_16_28), .i_b(w_carry_16_26), .i_c(w_carry_16_24), .ow_sum(w_sum_17_19), .ow_c(w_carry_17_19));
wire w_sum_17_17, w_carry_17_17;
math_adder_carry_save CSA_17_17(.i_a(w_carry_16_22), .i_b(w_carry_16_20), .i_c(w_carry_16_18), .ow_sum(w_sum_17_17), .ow_c(w_carry_17_17));
wire w_sum_17_15, w_carry_17_15;
math_adder_carry_save CSA_17_15(.i_a(w_carry_16_16), .i_b(w_carry_16_14), .i_c(w_carry_16_12), .ow_sum(w_sum_17_15), .ow_c(w_carry_17_15));
wire w_sum_17_13, w_carry_17_13;
math_adder_carry_save CSA_17_13(.i_a(w_carry_16_10), .i_b(w_carry_16_8), .i_c(w_carry_16_6), .ow_sum(w_sum_17_13), .ow_c(w_carry_17_13));
wire w_sum_17_11, w_carry_17_11;
math_adder_carry_save CSA_17_11(.i_a(w_carry_16_4), .i_b(w_carry_16_2), .i_c(w_sum_17_29), .ow_sum(w_sum_17_11), .ow_c(w_carry_17_11));
wire w_sum_17_9, w_carry_17_9;
math_adder_carry_save CSA_17_9(.i_a(w_sum_17_27), .i_b(w_sum_17_25), .i_c(w_sum_17_23), .ow_sum(w_sum_17_9), .ow_c(w_carry_17_9));
wire w_sum_17_7, w_carry_17_7;
math_adder_carry_save CSA_17_7(.i_a(w_sum_17_21), .i_b(w_sum_17_19), .i_c(w_sum_17_17), .ow_sum(w_sum_17_7), .ow_c(w_carry_17_7));
wire w_sum_17_5, w_carry_17_5;
math_adder_carry_save CSA_17_5(.i_a(w_sum_17_15), .i_b(w_sum_17_13), .i_c(w_sum_17_11), .ow_sum(w_sum_17_5), .ow_c(w_carry_17_5));
wire w_sum_17_3, w_carry_17_3;
math_adder_carry_save CSA_17_3(.i_a(w_sum_17_9), .i_b(w_sum_17_7), .i_c(w_sum_17_5), .ow_sum(w_sum_17_3), .ow_c(w_carry_17_3));
wire w_sum_18_27, w_carry_18_27;
math_adder_carry_save CSA_18_27(.i_a(w_pp_3_15), .i_b(w_pp_4_14), .i_c(w_pp_5_13), .ow_sum(w_sum_18_27), .ow_c(w_carry_18_27));
wire w_sum_18_25, w_carry_18_25;
math_adder_carry_save CSA_18_25(.i_a(w_pp_6_12), .i_b(w_pp_7_11), .i_c(w_pp_8_10), .ow_sum(w_sum_18_25), .ow_c(w_carry_18_25));
wire w_sum_18_23, w_carry_18_23;
math_adder_carry_save CSA_18_23(.i_a(w_pp_9_9), .i_b(w_pp_10_8), .i_c(w_pp_11_7), .ow_sum(w_sum_18_23), .ow_c(w_carry_18_23));
wire w_sum_18_21, w_carry_18_21;
math_adder_carry_save CSA_18_21(.i_a(w_pp_12_6), .i_b(w_pp_13_5), .i_c(w_pp_14_4), .ow_sum(w_sum_18_21), .ow_c(w_carry_18_21));
wire w_sum_18_19, w_carry_18_19;
math_adder_carry_save CSA_18_19(.i_a(w_pp_15_3), .i_b(w_carry_17_29), .i_c(w_carry_17_27), .ow_sum(w_sum_18_19), .ow_c(w_carry_18_19));
wire w_sum_18_17, w_carry_18_17;
math_adder_carry_save CSA_18_17(.i_a(w_carry_17_25), .i_b(w_carry_17_23), .i_c(w_carry_17_21), .ow_sum(w_sum_18_17), .ow_c(w_carry_18_17));
wire w_sum_18_15, w_carry_18_15;
math_adder_carry_save CSA_18_15(.i_a(w_carry_17_19), .i_b(w_carry_17_17), .i_c(w_carry_17_15), .ow_sum(w_sum_18_15), .ow_c(w_carry_18_15));
wire w_sum_18_13, w_carry_18_13;
math_adder_carry_save CSA_18_13(.i_a(w_carry_17_13), .i_b(w_carry_17_11), .i_c(w_carry_17_9), .ow_sum(w_sum_18_13), .ow_c(w_carry_18_13));
wire w_sum_18_11, w_carry_18_11;
math_adder_carry_save CSA_18_11(.i_a(w_carry_17_7), .i_b(w_carry_17_5), .i_c(w_carry_17_3), .ow_sum(w_sum_18_11), .ow_c(w_carry_18_11));
wire w_sum_18_9, w_carry_18_9;
math_adder_carry_save CSA_18_9(.i_a(w_sum_18_27), .i_b(w_sum_18_25), .i_c(w_sum_18_23), .ow_sum(w_sum_18_9), .ow_c(w_carry_18_9));
wire w_sum_18_7, w_carry_18_7;
math_adder_carry_save CSA_18_7(.i_a(w_sum_18_21), .i_b(w_sum_18_19), .i_c(w_sum_18_17), .ow_sum(w_sum_18_7), .ow_c(w_carry_18_7));
wire w_sum_18_5, w_carry_18_5;
math_adder_carry_save CSA_18_5(.i_a(w_sum_18_15), .i_b(w_sum_18_13), .i_c(w_sum_18_11), .ow_sum(w_sum_18_5), .ow_c(w_carry_18_5));
wire w_sum_18_3, w_carry_18_3;
math_adder_carry_save CSA_18_3(.i_a(w_sum_18_9), .i_b(w_sum_18_7), .i_c(w_sum_18_5), .ow_sum(w_sum_18_3), .ow_c(w_carry_18_3));
wire w_sum_19_25, w_carry_19_25;
math_adder_carry_save CSA_19_25(.i_a(w_pp_4_15), .i_b(w_pp_5_14), .i_c(w_pp_6_13), .ow_sum(w_sum_19_25), .ow_c(w_carry_19_25));
wire w_sum_19_23, w_carry_19_23;
math_adder_carry_save CSA_19_23(.i_a(w_pp_7_12), .i_b(w_pp_8_11), .i_c(w_pp_9_10), .ow_sum(w_sum_19_23), .ow_c(w_carry_19_23));
wire w_sum_19_21, w_carry_19_21;
math_adder_carry_save CSA_19_21(.i_a(w_pp_10_9), .i_b(w_pp_11_8), .i_c(w_pp_12_7), .ow_sum(w_sum_19_21), .ow_c(w_carry_19_21));
wire w_sum_19_19, w_carry_19_19;
math_adder_carry_save CSA_19_19(.i_a(w_pp_13_6), .i_b(w_pp_14_5), .i_c(w_pp_15_4), .ow_sum(w_sum_19_19), .ow_c(w_carry_19_19));
wire w_sum_19_17, w_carry_19_17;
math_adder_carry_save CSA_19_17(.i_a(w_carry_18_27), .i_b(w_carry_18_25), .i_c(w_carry_18_23), .ow_sum(w_sum_19_17), .ow_c(w_carry_19_17));
wire w_sum_19_15, w_carry_19_15;
math_adder_carry_save CSA_19_15(.i_a(w_carry_18_21), .i_b(w_carry_18_19), .i_c(w_carry_18_17), .ow_sum(w_sum_19_15), .ow_c(w_carry_19_15));
wire w_sum_19_13, w_carry_19_13;
math_adder_carry_save CSA_19_13(.i_a(w_carry_18_15), .i_b(w_carry_18_13), .i_c(w_carry_18_11), .ow_sum(w_sum_19_13), .ow_c(w_carry_19_13));
wire w_sum_19_11, w_carry_19_11;
math_adder_carry_save CSA_19_11(.i_a(w_carry_18_9), .i_b(w_carry_18_7), .i_c(w_carry_18_5), .ow_sum(w_sum_19_11), .ow_c(w_carry_19_11));
wire w_sum_19_9, w_carry_19_9;
math_adder_carry_save CSA_19_9(.i_a(w_carry_18_3), .i_b(w_sum_19_25), .i_c(w_sum_19_23), .ow_sum(w_sum_19_9), .ow_c(w_carry_19_9));
wire w_sum_19_7, w_carry_19_7;
math_adder_carry_save CSA_19_7(.i_a(w_sum_19_21), .i_b(w_sum_19_19), .i_c(w_sum_19_17), .ow_sum(w_sum_19_7), .ow_c(w_carry_19_7));
wire w_sum_19_5, w_carry_19_5;
math_adder_carry_save CSA_19_5(.i_a(w_sum_19_15), .i_b(w_sum_19_13), .i_c(w_sum_19_11), .ow_sum(w_sum_19_5), .ow_c(w_carry_19_5));
wire w_sum_19_3, w_carry_19_3;
math_adder_carry_save CSA_19_3(.i_a(w_sum_19_9), .i_b(w_sum_19_7), .i_c(w_sum_19_5), .ow_sum(w_sum_19_3), .ow_c(w_carry_19_3));
wire w_sum_20_23, w_carry_20_23;
math_adder_carry_save CSA_20_23(.i_a(w_pp_5_15), .i_b(w_pp_6_14), .i_c(w_pp_7_13), .ow_sum(w_sum_20_23), .ow_c(w_carry_20_23));
wire w_sum_20_21, w_carry_20_21;
math_adder_carry_save CSA_20_21(.i_a(w_pp_8_12), .i_b(w_pp_9_11), .i_c(w_pp_10_10), .ow_sum(w_sum_20_21), .ow_c(w_carry_20_21));
wire w_sum_20_19, w_carry_20_19;
math_adder_carry_save CSA_20_19(.i_a(w_pp_11_9), .i_b(w_pp_12_8), .i_c(w_pp_13_7), .ow_sum(w_sum_20_19), .ow_c(w_carry_20_19));
wire w_sum_20_17, w_carry_20_17;
math_adder_carry_save CSA_20_17(.i_a(w_pp_14_6), .i_b(w_pp_15_5), .i_c(w_carry_19_25), .ow_sum(w_sum_20_17), .ow_c(w_carry_20_17));
wire w_sum_20_15, w_carry_20_15;
math_adder_carry_save CSA_20_15(.i_a(w_carry_19_23), .i_b(w_carry_19_21), .i_c(w_carry_19_19), .ow_sum(w_sum_20_15), .ow_c(w_carry_20_15));
wire w_sum_20_13, w_carry_20_13;
math_adder_carry_save CSA_20_13(.i_a(w_carry_19_17), .i_b(w_carry_19_15), .i_c(w_carry_19_13), .ow_sum(w_sum_20_13), .ow_c(w_carry_20_13));
wire w_sum_20_11, w_carry_20_11;
math_adder_carry_save CSA_20_11(.i_a(w_carry_19_11), .i_b(w_carry_19_9), .i_c(w_carry_19_7), .ow_sum(w_sum_20_11), .ow_c(w_carry_20_11));
wire w_sum_20_9, w_carry_20_9;
math_adder_carry_save CSA_20_9(.i_a(w_carry_19_5), .i_b(w_carry_19_3), .i_c(w_sum_20_23), .ow_sum(w_sum_20_9), .ow_c(w_carry_20_9));
wire w_sum_20_7, w_carry_20_7;
math_adder_carry_save CSA_20_7(.i_a(w_sum_20_21), .i_b(w_sum_20_19), .i_c(w_sum_20_17), .ow_sum(w_sum_20_7), .ow_c(w_carry_20_7));
wire w_sum_20_5, w_carry_20_5;
math_adder_carry_save CSA_20_5(.i_a(w_sum_20_15), .i_b(w_sum_20_13), .i_c(w_sum_20_11), .ow_sum(w_sum_20_5), .ow_c(w_carry_20_5));
wire w_sum_20_3, w_carry_20_3;
math_adder_carry_save CSA_20_3(.i_a(w_sum_20_9), .i_b(w_sum_20_7), .i_c(w_sum_20_5), .ow_sum(w_sum_20_3), .ow_c(w_carry_20_3));
wire w_sum_21_21, w_carry_21_21;
math_adder_carry_save CSA_21_21(.i_a(w_pp_6_15), .i_b(w_pp_7_14), .i_c(w_pp_8_13), .ow_sum(w_sum_21_21), .ow_c(w_carry_21_21));
wire w_sum_21_19, w_carry_21_19;
math_adder_carry_save CSA_21_19(.i_a(w_pp_9_12), .i_b(w_pp_10_11), .i_c(w_pp_11_10), .ow_sum(w_sum_21_19), .ow_c(w_carry_21_19));
wire w_sum_21_17, w_carry_21_17;
math_adder_carry_save CSA_21_17(.i_a(w_pp_12_9), .i_b(w_pp_13_8), .i_c(w_pp_14_7), .ow_sum(w_sum_21_17), .ow_c(w_carry_21_17));
wire w_sum_21_15, w_carry_21_15;
math_adder_carry_save CSA_21_15(.i_a(w_pp_15_6), .i_b(w_carry_20_23), .i_c(w_carry_20_21), .ow_sum(w_sum_21_15), .ow_c(w_carry_21_15));
wire w_sum_21_13, w_carry_21_13;
math_adder_carry_save CSA_21_13(.i_a(w_carry_20_19), .i_b(w_carry_20_17), .i_c(w_carry_20_15), .ow_sum(w_sum_21_13), .ow_c(w_carry_21_13));
wire w_sum_21_11, w_carry_21_11;
math_adder_carry_save CSA_21_11(.i_a(w_carry_20_13), .i_b(w_carry_20_11), .i_c(w_carry_20_9), .ow_sum(w_sum_21_11), .ow_c(w_carry_21_11));
wire w_sum_21_9, w_carry_21_9;
math_adder_carry_save CSA_21_9(.i_a(w_carry_20_7), .i_b(w_carry_20_5), .i_c(w_carry_20_3), .ow_sum(w_sum_21_9), .ow_c(w_carry_21_9));
wire w_sum_21_7, w_carry_21_7;
math_adder_carry_save CSA_21_7(.i_a(w_sum_21_21), .i_b(w_sum_21_19), .i_c(w_sum_21_17), .ow_sum(w_sum_21_7), .ow_c(w_carry_21_7));
wire w_sum_21_5, w_carry_21_5;
math_adder_carry_save CSA_21_5(.i_a(w_sum_21_15), .i_b(w_sum_21_13), .i_c(w_sum_21_11), .ow_sum(w_sum_21_5), .ow_c(w_carry_21_5));
wire w_sum_21_3, w_carry_21_3;
math_adder_carry_save CSA_21_3(.i_a(w_sum_21_9), .i_b(w_sum_21_7), .i_c(w_sum_21_5), .ow_sum(w_sum_21_3), .ow_c(w_carry_21_3));
wire w_sum_22_19, w_carry_22_19;
math_adder_carry_save CSA_22_19(.i_a(w_pp_7_15), .i_b(w_pp_8_14), .i_c(w_pp_9_13), .ow_sum(w_sum_22_19), .ow_c(w_carry_22_19));
wire w_sum_22_17, w_carry_22_17;
math_adder_carry_save CSA_22_17(.i_a(w_pp_10_12), .i_b(w_pp_11_11), .i_c(w_pp_12_10), .ow_sum(w_sum_22_17), .ow_c(w_carry_22_17));
wire w_sum_22_15, w_carry_22_15;
math_adder_carry_save CSA_22_15(.i_a(w_pp_13_9), .i_b(w_pp_14_8), .i_c(w_pp_15_7), .ow_sum(w_sum_22_15), .ow_c(w_carry_22_15));
wire w_sum_22_13, w_carry_22_13;
math_adder_carry_save CSA_22_13(.i_a(w_carry_21_21), .i_b(w_carry_21_19), .i_c(w_carry_21_17), .ow_sum(w_sum_22_13), .ow_c(w_carry_22_13));
wire w_sum_22_11, w_carry_22_11;
math_adder_carry_save CSA_22_11(.i_a(w_carry_21_15), .i_b(w_carry_21_13), .i_c(w_carry_21_11), .ow_sum(w_sum_22_11), .ow_c(w_carry_22_11));
wire w_sum_22_9, w_carry_22_9;
math_adder_carry_save CSA_22_9(.i_a(w_carry_21_9), .i_b(w_carry_21_7), .i_c(w_carry_21_5), .ow_sum(w_sum_22_9), .ow_c(w_carry_22_9));
wire w_sum_22_7, w_carry_22_7;
math_adder_carry_save CSA_22_7(.i_a(w_carry_21_3), .i_b(w_sum_22_19), .i_c(w_sum_22_17), .ow_sum(w_sum_22_7), .ow_c(w_carry_22_7));
wire w_sum_22_5, w_carry_22_5;
math_adder_carry_save CSA_22_5(.i_a(w_sum_22_15), .i_b(w_sum_22_13), .i_c(w_sum_22_11), .ow_sum(w_sum_22_5), .ow_c(w_carry_22_5));
wire w_sum_22_3, w_carry_22_3;
math_adder_carry_save CSA_22_3(.i_a(w_sum_22_9), .i_b(w_sum_22_7), .i_c(w_sum_22_5), .ow_sum(w_sum_22_3), .ow_c(w_carry_22_3));
wire w_sum_23_17, w_carry_23_17;
math_adder_carry_save CSA_23_17(.i_a(w_pp_8_15), .i_b(w_pp_9_14), .i_c(w_pp_10_13), .ow_sum(w_sum_23_17), .ow_c(w_carry_23_17));
wire w_sum_23_15, w_carry_23_15;
math_adder_carry_save CSA_23_15(.i_a(w_pp_11_12), .i_b(w_pp_12_11), .i_c(w_pp_13_10), .ow_sum(w_sum_23_15), .ow_c(w_carry_23_15));
wire w_sum_23_13, w_carry_23_13;
math_adder_carry_save CSA_23_13(.i_a(w_pp_14_9), .i_b(w_pp_15_8), .i_c(w_carry_22_19), .ow_sum(w_sum_23_13), .ow_c(w_carry_23_13));
wire w_sum_23_11, w_carry_23_11;
math_adder_carry_save CSA_23_11(.i_a(w_carry_22_17), .i_b(w_carry_22_15), .i_c(w_carry_22_13), .ow_sum(w_sum_23_11), .ow_c(w_carry_23_11));
wire w_sum_23_9, w_carry_23_9;
math_adder_carry_save CSA_23_9(.i_a(w_carry_22_11), .i_b(w_carry_22_9), .i_c(w_carry_22_7), .ow_sum(w_sum_23_9), .ow_c(w_carry_23_9));
wire w_sum_23_7, w_carry_23_7;
math_adder_carry_save CSA_23_7(.i_a(w_carry_22_5), .i_b(w_carry_22_3), .i_c(w_sum_23_17), .ow_sum(w_sum_23_7), .ow_c(w_carry_23_7));
wire w_sum_23_5, w_carry_23_5;
math_adder_carry_save CSA_23_5(.i_a(w_sum_23_15), .i_b(w_sum_23_13), .i_c(w_sum_23_11), .ow_sum(w_sum_23_5), .ow_c(w_carry_23_5));
wire w_sum_23_3, w_carry_23_3;
math_adder_carry_save CSA_23_3(.i_a(w_sum_23_9), .i_b(w_sum_23_7), .i_c(w_sum_23_5), .ow_sum(w_sum_23_3), .ow_c(w_carry_23_3));
wire w_sum_24_15, w_carry_24_15;
math_adder_carry_save CSA_24_15(.i_a(w_pp_9_15), .i_b(w_pp_10_14), .i_c(w_pp_11_13), .ow_sum(w_sum_24_15), .ow_c(w_carry_24_15));
wire w_sum_24_13, w_carry_24_13;
math_adder_carry_save CSA_24_13(.i_a(w_pp_12_12), .i_b(w_pp_13_11), .i_c(w_pp_14_10), .ow_sum(w_sum_24_13), .ow_c(w_carry_24_13));
wire w_sum_24_11, w_carry_24_11;
math_adder_carry_save CSA_24_11(.i_a(w_pp_15_9), .i_b(w_carry_23_17), .i_c(w_carry_23_15), .ow_sum(w_sum_24_11), .ow_c(w_carry_24_11));
wire w_sum_24_9, w_carry_24_9;
math_adder_carry_save CSA_24_9(.i_a(w_carry_23_13), .i_b(w_carry_23_11), .i_c(w_carry_23_9), .ow_sum(w_sum_24_9), .ow_c(w_carry_24_9));
wire w_sum_24_7, w_carry_24_7;
math_adder_carry_save CSA_24_7(.i_a(w_carry_23_7), .i_b(w_carry_23_5), .i_c(w_carry_23_3), .ow_sum(w_sum_24_7), .ow_c(w_carry_24_7));
wire w_sum_24_5, w_carry_24_5;
math_adder_carry_save CSA_24_5(.i_a(w_sum_24_15), .i_b(w_sum_24_13), .i_c(w_sum_24_11), .ow_sum(w_sum_24_5), .ow_c(w_carry_24_5));
wire w_sum_24_3, w_carry_24_3;
math_adder_carry_save CSA_24_3(.i_a(w_sum_24_9), .i_b(w_sum_24_7), .i_c(w_sum_24_5), .ow_sum(w_sum_24_3), .ow_c(w_carry_24_3));
wire w_sum_25_13, w_carry_25_13;
math_adder_carry_save CSA_25_13(.i_a(w_pp_10_15), .i_b(w_pp_11_14), .i_c(w_pp_12_13), .ow_sum(w_sum_25_13), .ow_c(w_carry_25_13));
wire w_sum_25_11, w_carry_25_11;
math_adder_carry_save CSA_25_11(.i_a(w_pp_13_12), .i_b(w_pp_14_11), .i_c(w_pp_15_10), .ow_sum(w_sum_25_11), .ow_c(w_carry_25_11));
wire w_sum_25_9, w_carry_25_9;
math_adder_carry_save CSA_25_9(.i_a(w_carry_24_15), .i_b(w_carry_24_13), .i_c(w_carry_24_11), .ow_sum(w_sum_25_9), .ow_c(w_carry_25_9));
wire w_sum_25_7, w_carry_25_7;
math_adder_carry_save CSA_25_7(.i_a(w_carry_24_9), .i_b(w_carry_24_7), .i_c(w_carry_24_5), .ow_sum(w_sum_25_7), .ow_c(w_carry_25_7));
wire w_sum_25_5, w_carry_25_5;
math_adder_carry_save CSA_25_5(.i_a(w_carry_24_3), .i_b(w_sum_25_13), .i_c(w_sum_25_11), .ow_sum(w_sum_25_5), .ow_c(w_carry_25_5));
wire w_sum_25_3, w_carry_25_3;
math_adder_carry_save CSA_25_3(.i_a(w_sum_25_9), .i_b(w_sum_25_7), .i_c(w_sum_25_5), .ow_sum(w_sum_25_3), .ow_c(w_carry_25_3));
wire w_sum_26_11, w_carry_26_11;
math_adder_carry_save CSA_26_11(.i_a(w_pp_11_15), .i_b(w_pp_12_14), .i_c(w_pp_13_13), .ow_sum(w_sum_26_11), .ow_c(w_carry_26_11));
wire w_sum_26_9, w_carry_26_9;
math_adder_carry_save CSA_26_9(.i_a(w_pp_14_12), .i_b(w_pp_15_11), .i_c(w_carry_25_13), .ow_sum(w_sum_26_9), .ow_c(w_carry_26_9));
wire w_sum_26_7, w_carry_26_7;
math_adder_carry_save CSA_26_7(.i_a(w_carry_25_11), .i_b(w_carry_25_9), .i_c(w_carry_25_7), .ow_sum(w_sum_26_7), .ow_c(w_carry_26_7));
wire w_sum_26_5, w_carry_26_5;
math_adder_carry_save CSA_26_5(.i_a(w_carry_25_5), .i_b(w_carry_25_3), .i_c(w_sum_26_11), .ow_sum(w_sum_26_5), .ow_c(w_carry_26_5));
wire w_sum_26_3, w_carry_26_3;
math_adder_carry_save CSA_26_3(.i_a(w_sum_26_9), .i_b(w_sum_26_7), .i_c(w_sum_26_5), .ow_sum(w_sum_26_3), .ow_c(w_carry_26_3));
wire w_sum_27_9, w_carry_27_9;
math_adder_carry_save CSA_27_9(.i_a(w_pp_12_15), .i_b(w_pp_13_14), .i_c(w_pp_14_13), .ow_sum(w_sum_27_9), .ow_c(w_carry_27_9));
wire w_sum_27_7, w_carry_27_7;
math_adder_carry_save CSA_27_7(.i_a(w_pp_15_12), .i_b(w_carry_26_11), .i_c(w_carry_26_9), .ow_sum(w_sum_27_7), .ow_c(w_carry_27_7));
wire w_sum_27_5, w_carry_27_5;
math_adder_carry_save CSA_27_5(.i_a(w_carry_26_7), .i_b(w_carry_26_5), .i_c(w_carry_26_3), .ow_sum(w_sum_27_5), .ow_c(w_carry_27_5));
wire w_sum_27_3, w_carry_27_3;
math_adder_carry_save CSA_27_3(.i_a(w_sum_27_9), .i_b(w_sum_27_7), .i_c(w_sum_27_5), .ow_sum(w_sum_27_3), .ow_c(w_carry_27_3));
wire w_sum_28_7, w_carry_28_7;
math_adder_carry_save CSA_28_7(.i_a(w_pp_13_15), .i_b(w_pp_14_14), .i_c(w_pp_15_13), .ow_sum(w_sum_28_7), .ow_c(w_carry_28_7));
wire w_sum_28_5, w_carry_28_5;
math_adder_carry_save CSA_28_5(.i_a(w_carry_27_9), .i_b(w_carry_27_7), .i_c(w_carry_27_5), .ow_sum(w_sum_28_5), .ow_c(w_carry_28_5));
wire w_sum_28_3, w_carry_28_3;
math_adder_carry_save CSA_28_3(.i_a(w_carry_27_3), .i_b(w_sum_28_7), .i_c(w_sum_28_5), .ow_sum(w_sum_28_3), .ow_c(w_carry_28_3));
wire w_sum_29_5, w_carry_29_5;
math_adder_carry_save CSA_29_5(.i_a(w_pp_14_15), .i_b(w_pp_15_14), .i_c(w_carry_28_7), .ow_sum(w_sum_29_5), .ow_c(w_carry_29_5));
wire w_sum_29_3, w_carry_29_3;
math_adder_carry_save CSA_29_3(.i_a(w_carry_28_5), .i_b(w_carry_28_3), .i_c(w_sum_29_5), .ow_sum(w_sum_29_3), .ow_c(w_carry_29_3));
wire w_sum_30_3, w_carry_30_3;
math_adder_carry_save CSA_30_3(.i_a(w_pp_15_15), .i_b(w_carry_29_5), .i_c(w_carry_29_3), .ow_sum(w_sum_30_3), .ow_c(w_carry_30_3));

// Final product assignment
assign ow_product[0] = w_pp_0_0;
assign ow_product[1] = w_sum_1_2;
assign ow_product[2] = w_sum_2_2;
assign ow_product[3] = w_sum_3_2;
assign ow_product[4] = w_sum_4_2;
assign ow_product[5] = w_sum_5_2;
assign ow_product[6] = w_sum_6_2;
assign ow_product[7] = w_sum_7_2;
assign ow_product[8] = w_sum_8_2;
assign ow_product[9] = w_sum_9_2;
assign ow_product[10] = w_sum_10_2;
assign ow_product[11] = w_sum_11_2;
assign ow_product[12] = w_sum_12_2;
assign ow_product[13] = w_sum_13_2;
assign ow_product[14] = w_sum_14_2;
assign ow_product[15] = w_sum_15_2;
assign ow_product[16] = w_sum_16_2;
assign ow_product[17] = w_sum_17_3;
assign ow_product[18] = w_sum_18_3;
assign ow_product[19] = w_sum_19_3;
assign ow_product[20] = w_sum_20_3;
assign ow_product[21] = w_sum_21_3;
assign ow_product[22] = w_sum_22_3;
assign ow_product[23] = w_sum_23_3;
assign ow_product[24] = w_sum_24_3;
assign ow_product[25] = w_sum_25_3;
assign ow_product[26] = w_sum_26_3;
assign ow_product[27] = w_sum_27_3;
assign ow_product[28] = w_sum_28_3;
assign ow_product[29] = w_sum_29_3;
assign ow_product[30] = w_sum_30_3;
assign ow_product[31] = w_carry_30_3;


    // Debug purposes
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_wallace_tree_csa_16);
    end
                
endmodule : math_multiplier_wallace_tree_csa_16
