
`timescale 1ns / 1ps

module apb_xbar_wrap (
    input  logic                 clk,
    input  logic                 rst_n,

    input  logic                 m0_apb_psel,
    input  logic                 m0_apb_penable,
    input  logic                 m0_apb_pwrite,
    input  logic [AW-1:0]        m0_apb_paddr,
    input  logic [DW:0]          m0_apb_pwdata,
    input  logic [SW:0]          m0_apb_pstrb,
    output logic                 m0_apb_pready,
    output logic [DW:0]          m0_apb_prdata,
    output logic                 m0_apb_pslverr,

    input  logic                 m1_apb_psel,
    input  logic                 m1_apb_penable,
    input  logic                 m1_apb_pwrite,
    input  logic [AW-1:0]        m1_apb_paddr,
    input  logic [DW:0]          m1_apb_pwdata,
    input  logic [SW:0]          m1_apb_pstrb,
    output logic                 m1_apb_pready,
    output logic [DW:0]          m1_apb_prdata,
    output logic                 m1_apb_pslverr,

    input  logic                 m2_apb_psel,
    input  logic                 m2_apb_penable,
    input  logic                 m2_apb_pwrite,
    input  logic [AW-1:0]        m2_apb_paddr,
    input  logic [DW:0]          m2_apb_pwdata,
    input  logic [SW:0]          m2_apb_pstrb,
    output logic                 m2_apb_pready,
    output logic [DW:0]          m2_apb_prdata,
    output logic                 m2_apb_pslverr,

    output logic                 s0_apb_psel,
    output logic                 s0_apb_penable,
    output logic                 s0_apb_pwrite,
    output logic [AW-1:0]        s0_apb_paddr,
    output logic [DW-1:0]        s0_apb_pwdata,
    output logic [SW-1:0]        s0_apb_pstrb,
    input  logic                 s0_apb_pready,
    input  logic [DW-1:0]        s0_apb_prdata,
    input  logic                 s0_apb_pslverr,

    output logic                 s1_apb_psel,
    output logic                 s1_apb_penable,
    output logic                 s1_apb_pwrite,
    output logic [AW-1:0]        s1_apb_paddr,
    output logic [DW-1:0]        s1_apb_pwdata,
    output logic [SW-1:0]        s1_apb_pstrb,
    input  logic                 s1_apb_pready,
    input  logic [DW-1:0]        s1_apb_prdata,
    input  logic                 s1_apb_pslverr,

    output logic                 s2_apb_psel,
    output logic                 s2_apb_penable,
    output logic                 s2_apb_pwrite,
    output logic [AW-1:0]        s2_apb_paddr,
    output logic [DW-1:0]        s2_apb_pwdata,
    output logic [SW-1:0]        s2_apb_pstrb,
    input  logic                 s2_apb_pready,
    input  logic [DW-1:0]        s2_apb_prdata,
    input  logic                 s2_apb_pslverr,

    output logic                 s3_apb_psel,
    output logic                 s3_apb_penable,
    output logic                 s3_apb_pwrite,
    output logic [AW-1:0]        s3_apb_paddr,
    output logic [DW-1:0]        s3_apb_pwdata,
    output logic [SW-1:0]        s3_apb_pstrb,
    input  logic                 s3_apb_pready,
    input  logic [DW-1:0]        s3_apb_prdata,
    input  logic                 s3_apb_pslverr,

    output logic                 s4_apb_psel,
    output logic                 s4_apb_penable,
    output logic                 s4_apb_pwrite,
    output logic [AW-1:0]        s4_apb_paddr,
    output logic [DW-1:0]        s4_apb_pwdata,
    output logic [SW-1:0]        s4_apb_pstrb,
    input  logic                 s4_apb_pready,
    input  logic [DW-1:0]        s4_apb_prdata,
    input  logic                 s4_apb_pslverr
);


    localparam int DW  = DATA_WIDTH;
    localparam int AW  = ADDR_WIDTH;
    localparam int SW  = STRB_WIDTH;


    apb_xbar #(
        .M(3),
        .S(5),
        .ADDR_WIDTH(32),
        .DATA_WIDTH(32),
        .STRB_WIDTH(4),
    ) apb_xbar_inst (
        .clk(clk),
        .rst_n(rst_n),
        .SLAVE_ENABLE({1, 1, 1, 1, 1}),
        .SLAVE_ADDR_BASE('{32'h0, 32'h1000, 32'h2000, 32'h3000, 32'h4000}),
        .SLAVE_ADDR_LIMIT('{32'hFFF, 32'h1FFF, 32'h2FFF, 32'h3FFF, 32'h4FFF}),
        .THRESHOLDS('{4'h4, 4'h4, 4'h4, 4'h4, 4'h4})

        .m_apb_psel[0]     (m0_apb_psel),
        .m_apb_penable[0]  (m0_apb_penable),
        .m_apb_pwrite[0]   (m0_apb_pwrite),
        .m_apb_paddr[0]    (m0_apb_paddr),
        .m_apb_pwdata[0]   (m0_apb_pwdata),
        .m_apb_pstrb[0]    (m0_apb_pstrb),
        .m_apb_pready[0]   (m0_apb_pready),
        .m_apb_prdata[0]   (m0_apb_prdata),
        .m_apb_pslverr[0]  (m0_apb_pslverr),

        .m_apb_psel[1]     (m1_apb_psel),
        .m_apb_penable[1]  (m1_apb_penable),
        .m_apb_pwrite[1]   (m1_apb_pwrite),
        .m_apb_paddr[1]    (m1_apb_paddr),
        .m_apb_pwdata[1]   (m1_apb_pwdata),
        .m_apb_pstrb[1]    (m1_apb_pstrb),
        .m_apb_pready[1]   (m1_apb_pready),
        .m_apb_prdata[1]   (m1_apb_prdata),
        .m_apb_pslverr[1]  (m1_apb_pslverr),

        .m_apb_psel[2]     (m2_apb_psel),
        .m_apb_penable[2]  (m2_apb_penable),
        .m_apb_pwrite[2]   (m2_apb_pwrite),
        .m_apb_paddr[2]    (m2_apb_paddr),
        .m_apb_pwdata[2]   (m2_apb_pwdata),
        .m_apb_pstrb[2]    (m2_apb_pstrb),
        .m_apb_pready[2]   (m2_apb_pready),
        .m_apb_prdata[2]   (m2_apb_prdata),
        .m_apb_pslverr[2]  (m2_apb_pslverr),

        .s_apb_psel[0]    (s0_apb_psel),
        .s_apb_penable[0] (s0_apb_penable),
        .s_apb_pwrite[0]  (s0_apb_pwrite),
        .s_apb_paddr[0]   (s0_apb_paddr),
        .s_apb_pwdata[0]  (s0_apb_pwdata),
        .s_apb_pstrb[0]   (s0_apb_pstrb),
        .s_apb_pready[0]  (s0_apb_pready),
        .s_apb_prdata[0]  (s0_apb_prdata),
        .s_apb_pslverr[0] (s0_apb_pslverr),

        .s_apb_psel[1]    (s1_apb_psel),
        .s_apb_penable[1] (s1_apb_penable),
        .s_apb_pwrite[1]  (s1_apb_pwrite),
        .s_apb_paddr[1]   (s1_apb_paddr),
        .s_apb_pwdata[1]  (s1_apb_pwdata),
        .s_apb_pstrb[1]   (s1_apb_pstrb),
        .s_apb_pready[1]  (s1_apb_pready),
        .s_apb_prdata[1]  (s1_apb_prdata),
        .s_apb_pslverr[1] (s1_apb_pslverr),

        .s_apb_psel[2]    (s2_apb_psel),
        .s_apb_penable[2] (s2_apb_penable),
        .s_apb_pwrite[2]  (s2_apb_pwrite),
        .s_apb_paddr[2]   (s2_apb_paddr),
        .s_apb_pwdata[2]  (s2_apb_pwdata),
        .s_apb_pstrb[2]   (s2_apb_pstrb),
        .s_apb_pready[2]  (s2_apb_pready),
        .s_apb_prdata[2]  (s2_apb_prdata),
        .s_apb_pslverr[2] (s2_apb_pslverr),

        .s_apb_psel[3]    (s3_apb_psel),
        .s_apb_penable[3] (s3_apb_penable),
        .s_apb_pwrite[3]  (s3_apb_pwrite),
        .s_apb_paddr[3]   (s3_apb_paddr),
        .s_apb_pwdata[3]  (s3_apb_pwdata),
        .s_apb_pstrb[3]   (s3_apb_pstrb),
        .s_apb_pready[3]  (s3_apb_pready),
        .s_apb_prdata[3]  (s3_apb_prdata),
        .s_apb_pslverr[3] (s3_apb_pslverr),

        .s_apb_psel[4]    (s4_apb_psel),
        .s_apb_penable[4] (s4_apb_penable),
        .s_apb_pwrite[4]  (s4_apb_pwrite),
        .s_apb_paddr[4]   (s4_apb_paddr),
        .s_apb_pwdata[4]  (s4_apb_pwdata),
        .s_apb_pstrb[4]   (s4_apb_pstrb),
        .s_apb_pready[4]  (s4_apb_pready),
        .s_apb_prdata[4]  (s4_apb_prdata),
        .s_apb_pslverr[4] (s4_apb_pslverr)
    );

endmodule : apb_xbar_wrap
