// SPDX-License-Identifier: MIT
// SPDX-FileCopyrightText: 2024-2025 sean galloway
//
// RTL Design Sherpa - Industry-Standard RTL Design and Verification
// https://github.com/sean-galloway/RTLDesignSherpa
//
// Module: math_ieee754_2008_fp32_mantissa_mult
// Purpose: IEEE 754-2008 FP32 mantissa multiplier (24x24 with normalization and rounding)
//
// Documentation: IEEE754_ARCHITECTURE.md
// Subsystem: common
//
// Author: sean galloway
// Created: 2026-01-03
//
// AUTO-GENERATED FILE - DO NOT EDIT MANUALLY
// Generator: bin/rtl_generators/ieee754/fp32_mantissa_mult.py
// Regenerate: PYTHONPATH=bin:$PYTHONPATH python3 bin/rtl_generators/ieee754/generate_all.py rtl/common
//

`timescale 1ns / 1ps

module math_ieee754_2008_fp32_mantissa_mult(
    input  logic [22:0] i_mant_a,
    input  logic [22:0] i_mant_b,
    input  logic        i_a_is_normal,
    input  logic        i_b_is_normal,
    output logic [47:0] ow_product,
    output logic        ow_needs_norm,
    output logic [22:0] ow_mant_out,
    output logic        ow_round_bit,
    output logic        ow_sticky_bit
);

// Extend mantissa with implied leading 1 for normalized numbers
wire [23:0] w_mant_a_ext = {i_a_is_normal, i_mant_a};
wire [23:0] w_mant_b_ext = {i_b_is_normal, i_mant_b};

// 24x24 unsigned multiply using Dadda tree with 4:2 compressors
math_multiplier_dadda_4to2_024 u_mult (
    .i_multiplier(w_mant_a_ext),
    .i_multiplicand(w_mant_b_ext),
    .ow_product(ow_product)
);

// Normalization detection
// Product is in range [0, 4) before normalization
// If MSB (bit 47) is set: product >= 2.0, needs right shift
assign ow_needs_norm = ow_product[47];

// Extract result mantissa
// If needs_norm: take bits [46:24] (after implied 1)
// If not: take bits [45:23] (no shift needed)

// Normalized case:     1x.xxxxxxx...xxxxxxx -> take [46:24]
// Non-normalized case: 01.xxxxxxx...xxxxxxx -> take [45:23]
assign ow_mant_out = ow_needs_norm ? ow_product[46:24] : ow_product[45:23];

// Rounding support (Round-to-Nearest-Even)
// 
// For RNE, we need:
//   - Guard bit (G): first bit after mantissa
//   - Round bit (R): second bit after mantissa
//   - Sticky bit (S): OR of all remaining bits
// 
// If needs_norm (product >= 2):
//   mantissa = [46:24], G = [23], R = [22], S = |[21:0]
// If not needs_norm (product < 2):
//   mantissa = [45:23], G = [22], R = [21], S = |[20:0]

wire w_guard_norm    = ow_product[23];
wire w_guard_nonorm  = ow_product[22];

wire w_round_norm    = ow_product[22];
wire w_round_nonorm  = ow_product[21];

wire w_sticky_norm   = |ow_product[21:0];
wire w_sticky_nonorm = |ow_product[20:0];

assign ow_round_bit  = ow_needs_norm ? w_round_norm  : w_round_nonorm;
assign ow_sticky_bit = ow_needs_norm ? 
    (w_guard_norm | w_sticky_norm) : (w_guard_nonorm | w_sticky_nonorm);

endmodule
