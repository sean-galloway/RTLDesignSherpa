`timescale 1ns / 1ps

module math_multiplier_wallace_tree_016 #(
    parameter int N = 16
) (
    input  logic [  N-1:0] i_multiplier,
    input  logic [  N-1:0] i_multiplicand,
    output logic [2*N-1:0] ow_product
);

    // Partial Products
    wire w_pp_00_00 = i_multiplier[0] & i_multiplicand[0];
    wire w_pp_00_01 = i_multiplier[0] & i_multiplicand[1];
    wire w_pp_00_02 = i_multiplier[0] & i_multiplicand[2];
    wire w_pp_00_03 = i_multiplier[0] & i_multiplicand[3];
    wire w_pp_00_04 = i_multiplier[0] & i_multiplicand[4];
    wire w_pp_00_05 = i_multiplier[0] & i_multiplicand[5];
    wire w_pp_00_06 = i_multiplier[0] & i_multiplicand[6];
    wire w_pp_00_07 = i_multiplier[0] & i_multiplicand[7];
    wire w_pp_00_08 = i_multiplier[0] & i_multiplicand[8];
    wire w_pp_00_09 = i_multiplier[0] & i_multiplicand[9];
    wire w_pp_00_10 = i_multiplier[0] & i_multiplicand[10];
    wire w_pp_00_11 = i_multiplier[0] & i_multiplicand[11];
    wire w_pp_00_12 = i_multiplier[0] & i_multiplicand[12];
    wire w_pp_00_13 = i_multiplier[0] & i_multiplicand[13];
    wire w_pp_00_14 = i_multiplier[0] & i_multiplicand[14];
    wire w_pp_00_15 = i_multiplier[0] & i_multiplicand[15];
    wire w_pp_01_00 = i_multiplier[1] & i_multiplicand[0];
    wire w_pp_01_01 = i_multiplier[1] & i_multiplicand[1];
    wire w_pp_01_02 = i_multiplier[1] & i_multiplicand[2];
    wire w_pp_01_03 = i_multiplier[1] & i_multiplicand[3];
    wire w_pp_01_04 = i_multiplier[1] & i_multiplicand[4];
    wire w_pp_01_05 = i_multiplier[1] & i_multiplicand[5];
    wire w_pp_01_06 = i_multiplier[1] & i_multiplicand[6];
    wire w_pp_01_07 = i_multiplier[1] & i_multiplicand[7];
    wire w_pp_01_08 = i_multiplier[1] & i_multiplicand[8];
    wire w_pp_01_09 = i_multiplier[1] & i_multiplicand[9];
    wire w_pp_01_10 = i_multiplier[1] & i_multiplicand[10];
    wire w_pp_01_11 = i_multiplier[1] & i_multiplicand[11];
    wire w_pp_01_12 = i_multiplier[1] & i_multiplicand[12];
    wire w_pp_01_13 = i_multiplier[1] & i_multiplicand[13];
    wire w_pp_01_14 = i_multiplier[1] & i_multiplicand[14];
    wire w_pp_01_15 = i_multiplier[1] & i_multiplicand[15];
    wire w_pp_02_00 = i_multiplier[2] & i_multiplicand[0];
    wire w_pp_02_01 = i_multiplier[2] & i_multiplicand[1];
    wire w_pp_02_02 = i_multiplier[2] & i_multiplicand[2];
    wire w_pp_02_03 = i_multiplier[2] & i_multiplicand[3];
    wire w_pp_02_04 = i_multiplier[2] & i_multiplicand[4];
    wire w_pp_02_05 = i_multiplier[2] & i_multiplicand[5];
    wire w_pp_02_06 = i_multiplier[2] & i_multiplicand[6];
    wire w_pp_02_07 = i_multiplier[2] & i_multiplicand[7];
    wire w_pp_02_08 = i_multiplier[2] & i_multiplicand[8];
    wire w_pp_02_09 = i_multiplier[2] & i_multiplicand[9];
    wire w_pp_02_10 = i_multiplier[2] & i_multiplicand[10];
    wire w_pp_02_11 = i_multiplier[2] & i_multiplicand[11];
    wire w_pp_02_12 = i_multiplier[2] & i_multiplicand[12];
    wire w_pp_02_13 = i_multiplier[2] & i_multiplicand[13];
    wire w_pp_02_14 = i_multiplier[2] & i_multiplicand[14];
    wire w_pp_02_15 = i_multiplier[2] & i_multiplicand[15];
    wire w_pp_03_00 = i_multiplier[3] & i_multiplicand[0];
    wire w_pp_03_01 = i_multiplier[3] & i_multiplicand[1];
    wire w_pp_03_02 = i_multiplier[3] & i_multiplicand[2];
    wire w_pp_03_03 = i_multiplier[3] & i_multiplicand[3];
    wire w_pp_03_04 = i_multiplier[3] & i_multiplicand[4];
    wire w_pp_03_05 = i_multiplier[3] & i_multiplicand[5];
    wire w_pp_03_06 = i_multiplier[3] & i_multiplicand[6];
    wire w_pp_03_07 = i_multiplier[3] & i_multiplicand[7];
    wire w_pp_03_08 = i_multiplier[3] & i_multiplicand[8];
    wire w_pp_03_09 = i_multiplier[3] & i_multiplicand[9];
    wire w_pp_03_10 = i_multiplier[3] & i_multiplicand[10];
    wire w_pp_03_11 = i_multiplier[3] & i_multiplicand[11];
    wire w_pp_03_12 = i_multiplier[3] & i_multiplicand[12];
    wire w_pp_03_13 = i_multiplier[3] & i_multiplicand[13];
    wire w_pp_03_14 = i_multiplier[3] & i_multiplicand[14];
    wire w_pp_03_15 = i_multiplier[3] & i_multiplicand[15];
    wire w_pp_04_00 = i_multiplier[4] & i_multiplicand[0];
    wire w_pp_04_01 = i_multiplier[4] & i_multiplicand[1];
    wire w_pp_04_02 = i_multiplier[4] & i_multiplicand[2];
    wire w_pp_04_03 = i_multiplier[4] & i_multiplicand[3];
    wire w_pp_04_04 = i_multiplier[4] & i_multiplicand[4];
    wire w_pp_04_05 = i_multiplier[4] & i_multiplicand[5];
    wire w_pp_04_06 = i_multiplier[4] & i_multiplicand[6];
    wire w_pp_04_07 = i_multiplier[4] & i_multiplicand[7];
    wire w_pp_04_08 = i_multiplier[4] & i_multiplicand[8];
    wire w_pp_04_09 = i_multiplier[4] & i_multiplicand[9];
    wire w_pp_04_10 = i_multiplier[4] & i_multiplicand[10];
    wire w_pp_04_11 = i_multiplier[4] & i_multiplicand[11];
    wire w_pp_04_12 = i_multiplier[4] & i_multiplicand[12];
    wire w_pp_04_13 = i_multiplier[4] & i_multiplicand[13];
    wire w_pp_04_14 = i_multiplier[4] & i_multiplicand[14];
    wire w_pp_04_15 = i_multiplier[4] & i_multiplicand[15];
    wire w_pp_05_00 = i_multiplier[5] & i_multiplicand[0];
    wire w_pp_05_01 = i_multiplier[5] & i_multiplicand[1];
    wire w_pp_05_02 = i_multiplier[5] & i_multiplicand[2];
    wire w_pp_05_03 = i_multiplier[5] & i_multiplicand[3];
    wire w_pp_05_04 = i_multiplier[5] & i_multiplicand[4];
    wire w_pp_05_05 = i_multiplier[5] & i_multiplicand[5];
    wire w_pp_05_06 = i_multiplier[5] & i_multiplicand[6];
    wire w_pp_05_07 = i_multiplier[5] & i_multiplicand[7];
    wire w_pp_05_08 = i_multiplier[5] & i_multiplicand[8];
    wire w_pp_05_09 = i_multiplier[5] & i_multiplicand[9];
    wire w_pp_05_10 = i_multiplier[5] & i_multiplicand[10];
    wire w_pp_05_11 = i_multiplier[5] & i_multiplicand[11];
    wire w_pp_05_12 = i_multiplier[5] & i_multiplicand[12];
    wire w_pp_05_13 = i_multiplier[5] & i_multiplicand[13];
    wire w_pp_05_14 = i_multiplier[5] & i_multiplicand[14];
    wire w_pp_05_15 = i_multiplier[5] & i_multiplicand[15];
    wire w_pp_06_00 = i_multiplier[6] & i_multiplicand[0];
    wire w_pp_06_01 = i_multiplier[6] & i_multiplicand[1];
    wire w_pp_06_02 = i_multiplier[6] & i_multiplicand[2];
    wire w_pp_06_03 = i_multiplier[6] & i_multiplicand[3];
    wire w_pp_06_04 = i_multiplier[6] & i_multiplicand[4];
    wire w_pp_06_05 = i_multiplier[6] & i_multiplicand[5];
    wire w_pp_06_06 = i_multiplier[6] & i_multiplicand[6];
    wire w_pp_06_07 = i_multiplier[6] & i_multiplicand[7];
    wire w_pp_06_08 = i_multiplier[6] & i_multiplicand[8];
    wire w_pp_06_09 = i_multiplier[6] & i_multiplicand[9];
    wire w_pp_06_10 = i_multiplier[6] & i_multiplicand[10];
    wire w_pp_06_11 = i_multiplier[6] & i_multiplicand[11];
    wire w_pp_06_12 = i_multiplier[6] & i_multiplicand[12];
    wire w_pp_06_13 = i_multiplier[6] & i_multiplicand[13];
    wire w_pp_06_14 = i_multiplier[6] & i_multiplicand[14];
    wire w_pp_06_15 = i_multiplier[6] & i_multiplicand[15];
    wire w_pp_07_00 = i_multiplier[7] & i_multiplicand[0];
    wire w_pp_07_01 = i_multiplier[7] & i_multiplicand[1];
    wire w_pp_07_02 = i_multiplier[7] & i_multiplicand[2];
    wire w_pp_07_03 = i_multiplier[7] & i_multiplicand[3];
    wire w_pp_07_04 = i_multiplier[7] & i_multiplicand[4];
    wire w_pp_07_05 = i_multiplier[7] & i_multiplicand[5];
    wire w_pp_07_06 = i_multiplier[7] & i_multiplicand[6];
    wire w_pp_07_07 = i_multiplier[7] & i_multiplicand[7];
    wire w_pp_07_08 = i_multiplier[7] & i_multiplicand[8];
    wire w_pp_07_09 = i_multiplier[7] & i_multiplicand[9];
    wire w_pp_07_10 = i_multiplier[7] & i_multiplicand[10];
    wire w_pp_07_11 = i_multiplier[7] & i_multiplicand[11];
    wire w_pp_07_12 = i_multiplier[7] & i_multiplicand[12];
    wire w_pp_07_13 = i_multiplier[7] & i_multiplicand[13];
    wire w_pp_07_14 = i_multiplier[7] & i_multiplicand[14];
    wire w_pp_07_15 = i_multiplier[7] & i_multiplicand[15];
    wire w_pp_08_00 = i_multiplier[8] & i_multiplicand[0];
    wire w_pp_08_01 = i_multiplier[8] & i_multiplicand[1];
    wire w_pp_08_02 = i_multiplier[8] & i_multiplicand[2];
    wire w_pp_08_03 = i_multiplier[8] & i_multiplicand[3];
    wire w_pp_08_04 = i_multiplier[8] & i_multiplicand[4];
    wire w_pp_08_05 = i_multiplier[8] & i_multiplicand[5];
    wire w_pp_08_06 = i_multiplier[8] & i_multiplicand[6];
    wire w_pp_08_07 = i_multiplier[8] & i_multiplicand[7];
    wire w_pp_08_08 = i_multiplier[8] & i_multiplicand[8];
    wire w_pp_08_09 = i_multiplier[8] & i_multiplicand[9];
    wire w_pp_08_10 = i_multiplier[8] & i_multiplicand[10];
    wire w_pp_08_11 = i_multiplier[8] & i_multiplicand[11];
    wire w_pp_08_12 = i_multiplier[8] & i_multiplicand[12];
    wire w_pp_08_13 = i_multiplier[8] & i_multiplicand[13];
    wire w_pp_08_14 = i_multiplier[8] & i_multiplicand[14];
    wire w_pp_08_15 = i_multiplier[8] & i_multiplicand[15];
    wire w_pp_09_00 = i_multiplier[9] & i_multiplicand[0];
    wire w_pp_09_01 = i_multiplier[9] & i_multiplicand[1];
    wire w_pp_09_02 = i_multiplier[9] & i_multiplicand[2];
    wire w_pp_09_03 = i_multiplier[9] & i_multiplicand[3];
    wire w_pp_09_04 = i_multiplier[9] & i_multiplicand[4];
    wire w_pp_09_05 = i_multiplier[9] & i_multiplicand[5];
    wire w_pp_09_06 = i_multiplier[9] & i_multiplicand[6];
    wire w_pp_09_07 = i_multiplier[9] & i_multiplicand[7];
    wire w_pp_09_08 = i_multiplier[9] & i_multiplicand[8];
    wire w_pp_09_09 = i_multiplier[9] & i_multiplicand[9];
    wire w_pp_09_10 = i_multiplier[9] & i_multiplicand[10];
    wire w_pp_09_11 = i_multiplier[9] & i_multiplicand[11];
    wire w_pp_09_12 = i_multiplier[9] & i_multiplicand[12];
    wire w_pp_09_13 = i_multiplier[9] & i_multiplicand[13];
    wire w_pp_09_14 = i_multiplier[9] & i_multiplicand[14];
    wire w_pp_09_15 = i_multiplier[9] & i_multiplicand[15];
    wire w_pp_10_00 = i_multiplier[10] & i_multiplicand[0];
    wire w_pp_10_01 = i_multiplier[10] & i_multiplicand[1];
    wire w_pp_10_02 = i_multiplier[10] & i_multiplicand[2];
    wire w_pp_10_03 = i_multiplier[10] & i_multiplicand[3];
    wire w_pp_10_04 = i_multiplier[10] & i_multiplicand[4];
    wire w_pp_10_05 = i_multiplier[10] & i_multiplicand[5];
    wire w_pp_10_06 = i_multiplier[10] & i_multiplicand[6];
    wire w_pp_10_07 = i_multiplier[10] & i_multiplicand[7];
    wire w_pp_10_08 = i_multiplier[10] & i_multiplicand[8];
    wire w_pp_10_09 = i_multiplier[10] & i_multiplicand[9];
    wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
    wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
    wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
    wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
    wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
    wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
    wire w_pp_11_00 = i_multiplier[11] & i_multiplicand[0];
    wire w_pp_11_01 = i_multiplier[11] & i_multiplicand[1];
    wire w_pp_11_02 = i_multiplier[11] & i_multiplicand[2];
    wire w_pp_11_03 = i_multiplier[11] & i_multiplicand[3];
    wire w_pp_11_04 = i_multiplier[11] & i_multiplicand[4];
    wire w_pp_11_05 = i_multiplier[11] & i_multiplicand[5];
    wire w_pp_11_06 = i_multiplier[11] & i_multiplicand[6];
    wire w_pp_11_07 = i_multiplier[11] & i_multiplicand[7];
    wire w_pp_11_08 = i_multiplier[11] & i_multiplicand[8];
    wire w_pp_11_09 = i_multiplier[11] & i_multiplicand[9];
    wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
    wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
    wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
    wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
    wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
    wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
    wire w_pp_12_00 = i_multiplier[12] & i_multiplicand[0];
    wire w_pp_12_01 = i_multiplier[12] & i_multiplicand[1];
    wire w_pp_12_02 = i_multiplier[12] & i_multiplicand[2];
    wire w_pp_12_03 = i_multiplier[12] & i_multiplicand[3];
    wire w_pp_12_04 = i_multiplier[12] & i_multiplicand[4];
    wire w_pp_12_05 = i_multiplier[12] & i_multiplicand[5];
    wire w_pp_12_06 = i_multiplier[12] & i_multiplicand[6];
    wire w_pp_12_07 = i_multiplier[12] & i_multiplicand[7];
    wire w_pp_12_08 = i_multiplier[12] & i_multiplicand[8];
    wire w_pp_12_09 = i_multiplier[12] & i_multiplicand[9];
    wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
    wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
    wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
    wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
    wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
    wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
    wire w_pp_13_00 = i_multiplier[13] & i_multiplicand[0];
    wire w_pp_13_01 = i_multiplier[13] & i_multiplicand[1];
    wire w_pp_13_02 = i_multiplier[13] & i_multiplicand[2];
    wire w_pp_13_03 = i_multiplier[13] & i_multiplicand[3];
    wire w_pp_13_04 = i_multiplier[13] & i_multiplicand[4];
    wire w_pp_13_05 = i_multiplier[13] & i_multiplicand[5];
    wire w_pp_13_06 = i_multiplier[13] & i_multiplicand[6];
    wire w_pp_13_07 = i_multiplier[13] & i_multiplicand[7];
    wire w_pp_13_08 = i_multiplier[13] & i_multiplicand[8];
    wire w_pp_13_09 = i_multiplier[13] & i_multiplicand[9];
    wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
    wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
    wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
    wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
    wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
    wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
    wire w_pp_14_00 = i_multiplier[14] & i_multiplicand[0];
    wire w_pp_14_01 = i_multiplier[14] & i_multiplicand[1];
    wire w_pp_14_02 = i_multiplier[14] & i_multiplicand[2];
    wire w_pp_14_03 = i_multiplier[14] & i_multiplicand[3];
    wire w_pp_14_04 = i_multiplier[14] & i_multiplicand[4];
    wire w_pp_14_05 = i_multiplier[14] & i_multiplicand[5];
    wire w_pp_14_06 = i_multiplier[14] & i_multiplicand[6];
    wire w_pp_14_07 = i_multiplier[14] & i_multiplicand[7];
    wire w_pp_14_08 = i_multiplier[14] & i_multiplicand[8];
    wire w_pp_14_09 = i_multiplier[14] & i_multiplicand[9];
    wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
    wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
    wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
    wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
    wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
    wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
    wire w_pp_15_00 = i_multiplier[15] & i_multiplicand[0];
    wire w_pp_15_01 = i_multiplier[15] & i_multiplicand[1];
    wire w_pp_15_02 = i_multiplier[15] & i_multiplicand[2];
    wire w_pp_15_03 = i_multiplier[15] & i_multiplicand[3];
    wire w_pp_15_04 = i_multiplier[15] & i_multiplicand[4];
    wire w_pp_15_05 = i_multiplier[15] & i_multiplicand[5];
    wire w_pp_15_06 = i_multiplier[15] & i_multiplicand[6];
    wire w_pp_15_07 = i_multiplier[15] & i_multiplicand[7];
    wire w_pp_15_08 = i_multiplier[15] & i_multiplicand[8];
    wire w_pp_15_09 = i_multiplier[15] & i_multiplicand[9];
    wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
    wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
    wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
    wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
    wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
    wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];

    // Partial products reduction using Wallace tree
    wire w_sum_01_02, w_carry_01_02;
    math_adder_half HA_01_02 (
        .i_a(w_pp_00_01),
        .i_b(w_pp_01_00),
        .ow_sum(w_sum_01_02),
        .ow_carry(w_carry_01_02)
    );
    wire w_sum_02_04, w_carry_02_04;

    math_adder_full FA_02_04 (
        .i_a(w_pp_00_02),
        .i_b(w_pp_01_01),
        .i_c(w_pp_02_00),
        .ow_sum(w_sum_02_04),
        .ow_carry(w_carry_02_04)
    );
    wire w_sum_02_02, w_carry_02_02;
    math_adder_half HA_02_02 (
        .i_a(w_carry_01_02),
        .i_b(w_sum_02_04),
        .ow_sum(w_sum_02_02),
        .ow_carry(w_carry_02_02)
    );
    wire w_sum_03_06, w_carry_03_06;

    math_adder_full FA_03_06 (
        .i_a(w_pp_00_03),
        .i_b(w_pp_01_02),
        .i_c(w_pp_02_01),
        .ow_sum(w_sum_03_06),
        .ow_carry(w_carry_03_06)
    );
    wire w_sum_03_04, w_carry_03_04;

    math_adder_full FA_03_04 (
        .i_a(w_pp_03_00),
        .i_b(w_carry_02_04),
        .i_c(w_carry_02_02),
        .ow_sum(w_sum_03_04),
        .ow_carry(w_carry_03_04)
    );
    wire w_sum_03_02, w_carry_03_02;
    math_adder_half HA_03_02 (
        .i_a(w_sum_03_06),
        .i_b(w_sum_03_04),
        .ow_sum(w_sum_03_02),
        .ow_carry(w_carry_03_02)
    );
    wire w_sum_04_08, w_carry_04_08;

    math_adder_full FA_04_08 (
        .i_a(w_pp_00_04),
        .i_b(w_pp_01_03),
        .i_c(w_pp_02_02),
        .ow_sum(w_sum_04_08),
        .ow_carry(w_carry_04_08)
    );
    wire w_sum_04_06, w_carry_04_06;

    math_adder_full FA_04_06 (
        .i_a(w_pp_03_01),
        .i_b(w_pp_04_00),
        .i_c(w_carry_03_06),
        .ow_sum(w_sum_04_06),
        .ow_carry(w_carry_04_06)
    );
    wire w_sum_04_04, w_carry_04_04;

    math_adder_full FA_04_04 (
        .i_a(w_carry_03_04),
        .i_b(w_carry_03_02),
        .i_c(w_sum_04_08),
        .ow_sum(w_sum_04_04),
        .ow_carry(w_carry_04_04)
    );
    wire w_sum_04_02, w_carry_04_02;
    math_adder_half HA_04_02 (
        .i_a(w_sum_04_06),
        .i_b(w_sum_04_04),
        .ow_sum(w_sum_04_02),
        .ow_carry(w_carry_04_02)
    );
    wire w_sum_05_10, w_carry_05_10;

    math_adder_full FA_05_10 (
        .i_a(w_pp_00_05),
        .i_b(w_pp_01_04),
        .i_c(w_pp_02_03),
        .ow_sum(w_sum_05_10),
        .ow_carry(w_carry_05_10)
    );
    wire w_sum_05_08, w_carry_05_08;

    math_adder_full FA_05_08 (
        .i_a(w_pp_03_02),
        .i_b(w_pp_04_01),
        .i_c(w_pp_05_00),
        .ow_sum(w_sum_05_08),
        .ow_carry(w_carry_05_08)
    );
    wire w_sum_05_06, w_carry_05_06;

    math_adder_full FA_05_06 (
        .i_a(w_carry_04_08),
        .i_b(w_carry_04_06),
        .i_c(w_carry_04_04),
        .ow_sum(w_sum_05_06),
        .ow_carry(w_carry_05_06)
    );
    wire w_sum_05_04, w_carry_05_04;

    math_adder_full FA_05_04 (
        .i_a(w_carry_04_02),
        .i_b(w_sum_05_10),
        .i_c(w_sum_05_08),
        .ow_sum(w_sum_05_04),
        .ow_carry(w_carry_05_04)
    );
    wire w_sum_05_02, w_carry_05_02;
    math_adder_half HA_05_02 (
        .i_a(w_sum_05_06),
        .i_b(w_sum_05_04),
        .ow_sum(w_sum_05_02),
        .ow_carry(w_carry_05_02)
    );
    wire w_sum_06_12, w_carry_06_12;

    math_adder_full FA_06_12 (
        .i_a(w_pp_00_06),
        .i_b(w_pp_01_05),
        .i_c(w_pp_02_04),
        .ow_sum(w_sum_06_12),
        .ow_carry(w_carry_06_12)
    );
    wire w_sum_06_10, w_carry_06_10;

    math_adder_full FA_06_10 (
        .i_a(w_pp_03_03),
        .i_b(w_pp_04_02),
        .i_c(w_pp_05_01),
        .ow_sum(w_sum_06_10),
        .ow_carry(w_carry_06_10)
    );
    wire w_sum_06_08, w_carry_06_08;

    math_adder_full FA_06_08 (
        .i_a(w_pp_06_00),
        .i_b(w_carry_05_10),
        .i_c(w_carry_05_08),
        .ow_sum(w_sum_06_08),
        .ow_carry(w_carry_06_08)
    );
    wire w_sum_06_06, w_carry_06_06;

    math_adder_full FA_06_06 (
        .i_a(w_carry_05_06),
        .i_b(w_carry_05_04),
        .i_c(w_carry_05_02),
        .ow_sum(w_sum_06_06),
        .ow_carry(w_carry_06_06)
    );
    wire w_sum_06_04, w_carry_06_04;

    math_adder_full FA_06_04 (
        .i_a(w_sum_06_12),
        .i_b(w_sum_06_10),
        .i_c(w_sum_06_08),
        .ow_sum(w_sum_06_04),
        .ow_carry(w_carry_06_04)
    );
    wire w_sum_06_02, w_carry_06_02;
    math_adder_half HA_06_02 (
        .i_a(w_sum_06_06),
        .i_b(w_sum_06_04),
        .ow_sum(w_sum_06_02),
        .ow_carry(w_carry_06_02)
    );
    wire w_sum_07_14, w_carry_07_14;

    math_adder_full FA_07_14 (
        .i_a(w_pp_00_07),
        .i_b(w_pp_01_06),
        .i_c(w_pp_02_05),
        .ow_sum(w_sum_07_14),
        .ow_carry(w_carry_07_14)
    );
    wire w_sum_07_12, w_carry_07_12;

    math_adder_full FA_07_12 (
        .i_a(w_pp_03_04),
        .i_b(w_pp_04_03),
        .i_c(w_pp_05_02),
        .ow_sum(w_sum_07_12),
        .ow_carry(w_carry_07_12)
    );
    wire w_sum_07_10, w_carry_07_10;

    math_adder_full FA_07_10 (
        .i_a(w_pp_06_01),
        .i_b(w_pp_07_00),
        .i_c(w_carry_06_12),
        .ow_sum(w_sum_07_10),
        .ow_carry(w_carry_07_10)
    );
    wire w_sum_07_08, w_carry_07_08;

    math_adder_full FA_07_08 (
        .i_a(w_carry_06_10),
        .i_b(w_carry_06_08),
        .i_c(w_carry_06_06),
        .ow_sum(w_sum_07_08),
        .ow_carry(w_carry_07_08)
    );
    wire w_sum_07_06, w_carry_07_06;

    math_adder_full FA_07_06 (
        .i_a(w_carry_06_04),
        .i_b(w_carry_06_02),
        .i_c(w_sum_07_14),
        .ow_sum(w_sum_07_06),
        .ow_carry(w_carry_07_06)
    );
    wire w_sum_07_04, w_carry_07_04;

    math_adder_full FA_07_04 (
        .i_a(w_sum_07_12),
        .i_b(w_sum_07_10),
        .i_c(w_sum_07_08),
        .ow_sum(w_sum_07_04),
        .ow_carry(w_carry_07_04)
    );
    wire w_sum_07_02, w_carry_07_02;
    math_adder_half HA_07_02 (
        .i_a(w_sum_07_06),
        .i_b(w_sum_07_04),
        .ow_sum(w_sum_07_02),
        .ow_carry(w_carry_07_02)
    );
    wire w_sum_08_16, w_carry_08_16;

    math_adder_full FA_08_16 (
        .i_a(w_pp_00_08),
        .i_b(w_pp_01_07),
        .i_c(w_pp_02_06),
        .ow_sum(w_sum_08_16),
        .ow_carry(w_carry_08_16)
    );
    wire w_sum_08_14, w_carry_08_14;

    math_adder_full FA_08_14 (
        .i_a(w_pp_03_05),
        .i_b(w_pp_04_04),
        .i_c(w_pp_05_03),
        .ow_sum(w_sum_08_14),
        .ow_carry(w_carry_08_14)
    );
    wire w_sum_08_12, w_carry_08_12;

    math_adder_full FA_08_12 (
        .i_a(w_pp_06_02),
        .i_b(w_pp_07_01),
        .i_c(w_pp_08_00),
        .ow_sum(w_sum_08_12),
        .ow_carry(w_carry_08_12)
    );
    wire w_sum_08_10, w_carry_08_10;

    math_adder_full FA_08_10 (
        .i_a(w_carry_07_14),
        .i_b(w_carry_07_12),
        .i_c(w_carry_07_10),
        .ow_sum(w_sum_08_10),
        .ow_carry(w_carry_08_10)
    );
    wire w_sum_08_08, w_carry_08_08;

    math_adder_full FA_08_08 (
        .i_a(w_carry_07_08),
        .i_b(w_carry_07_06),
        .i_c(w_carry_07_04),
        .ow_sum(w_sum_08_08),
        .ow_carry(w_carry_08_08)
    );
    wire w_sum_08_06, w_carry_08_06;

    math_adder_full FA_08_06 (
        .i_a(w_carry_07_02),
        .i_b(w_sum_08_16),
        .i_c(w_sum_08_14),
        .ow_sum(w_sum_08_06),
        .ow_carry(w_carry_08_06)
    );
    wire w_sum_08_04, w_carry_08_04;

    math_adder_full FA_08_04 (
        .i_a(w_sum_08_12),
        .i_b(w_sum_08_10),
        .i_c(w_sum_08_08),
        .ow_sum(w_sum_08_04),
        .ow_carry(w_carry_08_04)
    );
    wire w_sum_08_02, w_carry_08_02;
    math_adder_half HA_08_02 (
        .i_a(w_sum_08_06),
        .i_b(w_sum_08_04),
        .ow_sum(w_sum_08_02),
        .ow_carry(w_carry_08_02)
    );
    wire w_sum_09_18, w_carry_09_18;

    math_adder_full FA_09_18 (
        .i_a(w_pp_00_09),
        .i_b(w_pp_01_08),
        .i_c(w_pp_02_07),
        .ow_sum(w_sum_09_18),
        .ow_carry(w_carry_09_18)
    );
    wire w_sum_09_16, w_carry_09_16;

    math_adder_full FA_09_16 (
        .i_a(w_pp_03_06),
        .i_b(w_pp_04_05),
        .i_c(w_pp_05_04),
        .ow_sum(w_sum_09_16),
        .ow_carry(w_carry_09_16)
    );
    wire w_sum_09_14, w_carry_09_14;

    math_adder_full FA_09_14 (
        .i_a(w_pp_06_03),
        .i_b(w_pp_07_02),
        .i_c(w_pp_08_01),
        .ow_sum(w_sum_09_14),
        .ow_carry(w_carry_09_14)
    );
    wire w_sum_09_12, w_carry_09_12;

    math_adder_full FA_09_12 (
        .i_a(w_pp_09_00),
        .i_b(w_carry_08_16),
        .i_c(w_carry_08_14),
        .ow_sum(w_sum_09_12),
        .ow_carry(w_carry_09_12)
    );
    wire w_sum_09_10, w_carry_09_10;

    math_adder_full FA_09_10 (
        .i_a(w_carry_08_12),
        .i_b(w_carry_08_10),
        .i_c(w_carry_08_08),
        .ow_sum(w_sum_09_10),
        .ow_carry(w_carry_09_10)
    );
    wire w_sum_09_08, w_carry_09_08;

    math_adder_full FA_09_08 (
        .i_a(w_carry_08_06),
        .i_b(w_carry_08_04),
        .i_c(w_carry_08_02),
        .ow_sum(w_sum_09_08),
        .ow_carry(w_carry_09_08)
    );
    wire w_sum_09_06, w_carry_09_06;

    math_adder_full FA_09_06 (
        .i_a(w_sum_09_18),
        .i_b(w_sum_09_16),
        .i_c(w_sum_09_14),
        .ow_sum(w_sum_09_06),
        .ow_carry(w_carry_09_06)
    );
    wire w_sum_09_04, w_carry_09_04;

    math_adder_full FA_09_04 (
        .i_a(w_sum_09_12),
        .i_b(w_sum_09_10),
        .i_c(w_sum_09_08),
        .ow_sum(w_sum_09_04),
        .ow_carry(w_carry_09_04)
    );
    wire w_sum_09_02, w_carry_09_02;
    math_adder_half HA_09_02 (
        .i_a(w_sum_09_06),
        .i_b(w_sum_09_04),
        .ow_sum(w_sum_09_02),
        .ow_carry(w_carry_09_02)
    );
    wire w_sum_10_20, w_carry_10_20;

    math_adder_full FA_10_20 (
        .i_a(w_pp_00_10),
        .i_b(w_pp_01_09),
        .i_c(w_pp_02_08),
        .ow_sum(w_sum_10_20),
        .ow_carry(w_carry_10_20)
    );
    wire w_sum_10_18, w_carry_10_18;

    math_adder_full FA_10_18 (
        .i_a(w_pp_03_07),
        .i_b(w_pp_04_06),
        .i_c(w_pp_05_05),
        .ow_sum(w_sum_10_18),
        .ow_carry(w_carry_10_18)
    );
    wire w_sum_10_16, w_carry_10_16;

    math_adder_full FA_10_16 (
        .i_a(w_pp_06_04),
        .i_b(w_pp_07_03),
        .i_c(w_pp_08_02),
        .ow_sum(w_sum_10_16),
        .ow_carry(w_carry_10_16)
    );
    wire w_sum_10_14, w_carry_10_14;

    math_adder_full FA_10_14 (
        .i_a(w_pp_09_01),
        .i_b(w_pp_10_00),
        .i_c(w_carry_09_18),
        .ow_sum(w_sum_10_14),
        .ow_carry(w_carry_10_14)
    );
    wire w_sum_10_12, w_carry_10_12;

    math_adder_full FA_10_12 (
        .i_a(w_carry_09_16),
        .i_b(w_carry_09_14),
        .i_c(w_carry_09_12),
        .ow_sum(w_sum_10_12),
        .ow_carry(w_carry_10_12)
    );
    wire w_sum_10_10, w_carry_10_10;

    math_adder_full FA_10_10 (
        .i_a(w_carry_09_10),
        .i_b(w_carry_09_08),
        .i_c(w_carry_09_06),
        .ow_sum(w_sum_10_10),
        .ow_carry(w_carry_10_10)
    );
    wire w_sum_10_08, w_carry_10_08;

    math_adder_full FA_10_08 (
        .i_a(w_carry_09_04),
        .i_b(w_carry_09_02),
        .i_c(w_sum_10_20),
        .ow_sum(w_sum_10_08),
        .ow_carry(w_carry_10_08)
    );
    wire w_sum_10_06, w_carry_10_06;

    math_adder_full FA_10_06 (
        .i_a(w_sum_10_18),
        .i_b(w_sum_10_16),
        .i_c(w_sum_10_14),
        .ow_sum(w_sum_10_06),
        .ow_carry(w_carry_10_06)
    );
    wire w_sum_10_04, w_carry_10_04;

    math_adder_full FA_10_04 (
        .i_a(w_sum_10_12),
        .i_b(w_sum_10_10),
        .i_c(w_sum_10_08),
        .ow_sum(w_sum_10_04),
        .ow_carry(w_carry_10_04)
    );
    wire w_sum_10_02, w_carry_10_02;
    math_adder_half HA_10_02 (
        .i_a(w_sum_10_06),
        .i_b(w_sum_10_04),
        .ow_sum(w_sum_10_02),
        .ow_carry(w_carry_10_02)
    );
    wire w_sum_11_22, w_carry_11_22;

    math_adder_full FA_11_22 (
        .i_a(w_pp_00_11),
        .i_b(w_pp_01_10),
        .i_c(w_pp_02_09),
        .ow_sum(w_sum_11_22),
        .ow_carry(w_carry_11_22)
    );
    wire w_sum_11_20, w_carry_11_20;

    math_adder_full FA_11_20 (
        .i_a(w_pp_03_08),
        .i_b(w_pp_04_07),
        .i_c(w_pp_05_06),
        .ow_sum(w_sum_11_20),
        .ow_carry(w_carry_11_20)
    );
    wire w_sum_11_18, w_carry_11_18;

    math_adder_full FA_11_18 (
        .i_a(w_pp_06_05),
        .i_b(w_pp_07_04),
        .i_c(w_pp_08_03),
        .ow_sum(w_sum_11_18),
        .ow_carry(w_carry_11_18)
    );
    wire w_sum_11_16, w_carry_11_16;

    math_adder_full FA_11_16 (
        .i_a(w_pp_09_02),
        .i_b(w_pp_10_01),
        .i_c(w_pp_11_00),
        .ow_sum(w_sum_11_16),
        .ow_carry(w_carry_11_16)
    );
    wire w_sum_11_14, w_carry_11_14;

    math_adder_full FA_11_14 (
        .i_a(w_carry_10_20),
        .i_b(w_carry_10_18),
        .i_c(w_carry_10_16),
        .ow_sum(w_sum_11_14),
        .ow_carry(w_carry_11_14)
    );
    wire w_sum_11_12, w_carry_11_12;

    math_adder_full FA_11_12 (
        .i_a(w_carry_10_14),
        .i_b(w_carry_10_12),
        .i_c(w_carry_10_10),
        .ow_sum(w_sum_11_12),
        .ow_carry(w_carry_11_12)
    );
    wire w_sum_11_10, w_carry_11_10;

    math_adder_full FA_11_10 (
        .i_a(w_carry_10_08),
        .i_b(w_carry_10_06),
        .i_c(w_carry_10_04),
        .ow_sum(w_sum_11_10),
        .ow_carry(w_carry_11_10)
    );
    wire w_sum_11_08, w_carry_11_08;

    math_adder_full FA_11_08 (
        .i_a(w_carry_10_02),
        .i_b(w_sum_11_22),
        .i_c(w_sum_11_20),
        .ow_sum(w_sum_11_08),
        .ow_carry(w_carry_11_08)
    );
    wire w_sum_11_06, w_carry_11_06;

    math_adder_full FA_11_06 (
        .i_a(w_sum_11_18),
        .i_b(w_sum_11_16),
        .i_c(w_sum_11_14),
        .ow_sum(w_sum_11_06),
        .ow_carry(w_carry_11_06)
    );
    wire w_sum_11_04, w_carry_11_04;

    math_adder_full FA_11_04 (
        .i_a(w_sum_11_12),
        .i_b(w_sum_11_10),
        .i_c(w_sum_11_08),
        .ow_sum(w_sum_11_04),
        .ow_carry(w_carry_11_04)
    );
    wire w_sum_11_02, w_carry_11_02;
    math_adder_half HA_11_02 (
        .i_a(w_sum_11_06),
        .i_b(w_sum_11_04),
        .ow_sum(w_sum_11_02),
        .ow_carry(w_carry_11_02)
    );
    wire w_sum_12_24, w_carry_12_24;

    math_adder_full FA_12_24 (
        .i_a(w_pp_00_12),
        .i_b(w_pp_01_11),
        .i_c(w_pp_02_10),
        .ow_sum(w_sum_12_24),
        .ow_carry(w_carry_12_24)
    );
    wire w_sum_12_22, w_carry_12_22;

    math_adder_full FA_12_22 (
        .i_a(w_pp_03_09),
        .i_b(w_pp_04_08),
        .i_c(w_pp_05_07),
        .ow_sum(w_sum_12_22),
        .ow_carry(w_carry_12_22)
    );
    wire w_sum_12_20, w_carry_12_20;

    math_adder_full FA_12_20 (
        .i_a(w_pp_06_06),
        .i_b(w_pp_07_05),
        .i_c(w_pp_08_04),
        .ow_sum(w_sum_12_20),
        .ow_carry(w_carry_12_20)
    );
    wire w_sum_12_18, w_carry_12_18;

    math_adder_full FA_12_18 (
        .i_a(w_pp_09_03),
        .i_b(w_pp_10_02),
        .i_c(w_pp_11_01),
        .ow_sum(w_sum_12_18),
        .ow_carry(w_carry_12_18)
    );
    wire w_sum_12_16, w_carry_12_16;

    math_adder_full FA_12_16 (
        .i_a(w_pp_12_00),
        .i_b(w_carry_11_22),
        .i_c(w_carry_11_20),
        .ow_sum(w_sum_12_16),
        .ow_carry(w_carry_12_16)
    );
    wire w_sum_12_14, w_carry_12_14;

    math_adder_full FA_12_14 (
        .i_a(w_carry_11_18),
        .i_b(w_carry_11_16),
        .i_c(w_carry_11_14),
        .ow_sum(w_sum_12_14),
        .ow_carry(w_carry_12_14)
    );
    wire w_sum_12_12, w_carry_12_12;

    math_adder_full FA_12_12 (
        .i_a(w_carry_11_12),
        .i_b(w_carry_11_10),
        .i_c(w_carry_11_08),
        .ow_sum(w_sum_12_12),
        .ow_carry(w_carry_12_12)
    );
    wire w_sum_12_10, w_carry_12_10;

    math_adder_full FA_12_10 (
        .i_a(w_carry_11_06),
        .i_b(w_carry_11_04),
        .i_c(w_carry_11_02),
        .ow_sum(w_sum_12_10),
        .ow_carry(w_carry_12_10)
    );
    wire w_sum_12_08, w_carry_12_08;

    math_adder_full FA_12_08 (
        .i_a(w_sum_12_24),
        .i_b(w_sum_12_22),
        .i_c(w_sum_12_20),
        .ow_sum(w_sum_12_08),
        .ow_carry(w_carry_12_08)
    );
    wire w_sum_12_06, w_carry_12_06;

    math_adder_full FA_12_06 (
        .i_a(w_sum_12_18),
        .i_b(w_sum_12_16),
        .i_c(w_sum_12_14),
        .ow_sum(w_sum_12_06),
        .ow_carry(w_carry_12_06)
    );
    wire w_sum_12_04, w_carry_12_04;

    math_adder_full FA_12_04 (
        .i_a(w_sum_12_12),
        .i_b(w_sum_12_10),
        .i_c(w_sum_12_08),
        .ow_sum(w_sum_12_04),
        .ow_carry(w_carry_12_04)
    );
    wire w_sum_12_02, w_carry_12_02;
    math_adder_half HA_12_02 (
        .i_a(w_sum_12_06),
        .i_b(w_sum_12_04),
        .ow_sum(w_sum_12_02),
        .ow_carry(w_carry_12_02)
    );
    wire w_sum_13_26, w_carry_13_26;

    math_adder_full FA_13_26 (
        .i_a(w_pp_00_13),
        .i_b(w_pp_01_12),
        .i_c(w_pp_02_11),
        .ow_sum(w_sum_13_26),
        .ow_carry(w_carry_13_26)
    );
    wire w_sum_13_24, w_carry_13_24;

    math_adder_full FA_13_24 (
        .i_a(w_pp_03_10),
        .i_b(w_pp_04_09),
        .i_c(w_pp_05_08),
        .ow_sum(w_sum_13_24),
        .ow_carry(w_carry_13_24)
    );
    wire w_sum_13_22, w_carry_13_22;

    math_adder_full FA_13_22 (
        .i_a(w_pp_06_07),
        .i_b(w_pp_07_06),
        .i_c(w_pp_08_05),
        .ow_sum(w_sum_13_22),
        .ow_carry(w_carry_13_22)
    );
    wire w_sum_13_20, w_carry_13_20;

    math_adder_full FA_13_20 (
        .i_a(w_pp_09_04),
        .i_b(w_pp_10_03),
        .i_c(w_pp_11_02),
        .ow_sum(w_sum_13_20),
        .ow_carry(w_carry_13_20)
    );
    wire w_sum_13_18, w_carry_13_18;

    math_adder_full FA_13_18 (
        .i_a(w_pp_12_01),
        .i_b(w_pp_13_00),
        .i_c(w_carry_12_24),
        .ow_sum(w_sum_13_18),
        .ow_carry(w_carry_13_18)
    );
    wire w_sum_13_16, w_carry_13_16;

    math_adder_full FA_13_16 (
        .i_a(w_carry_12_22),
        .i_b(w_carry_12_20),
        .i_c(w_carry_12_18),
        .ow_sum(w_sum_13_16),
        .ow_carry(w_carry_13_16)
    );
    wire w_sum_13_14, w_carry_13_14;

    math_adder_full FA_13_14 (
        .i_a(w_carry_12_16),
        .i_b(w_carry_12_14),
        .i_c(w_carry_12_12),
        .ow_sum(w_sum_13_14),
        .ow_carry(w_carry_13_14)
    );
    wire w_sum_13_12, w_carry_13_12;

    math_adder_full FA_13_12 (
        .i_a(w_carry_12_10),
        .i_b(w_carry_12_08),
        .i_c(w_carry_12_06),
        .ow_sum(w_sum_13_12),
        .ow_carry(w_carry_13_12)
    );
    wire w_sum_13_10, w_carry_13_10;

    math_adder_full FA_13_10 (
        .i_a(w_carry_12_04),
        .i_b(w_carry_12_02),
        .i_c(w_sum_13_26),
        .ow_sum(w_sum_13_10),
        .ow_carry(w_carry_13_10)
    );
    wire w_sum_13_08, w_carry_13_08;

    math_adder_full FA_13_08 (
        .i_a(w_sum_13_24),
        .i_b(w_sum_13_22),
        .i_c(w_sum_13_20),
        .ow_sum(w_sum_13_08),
        .ow_carry(w_carry_13_08)
    );
    wire w_sum_13_06, w_carry_13_06;

    math_adder_full FA_13_06 (
        .i_a(w_sum_13_18),
        .i_b(w_sum_13_16),
        .i_c(w_sum_13_14),
        .ow_sum(w_sum_13_06),
        .ow_carry(w_carry_13_06)
    );
    wire w_sum_13_04, w_carry_13_04;

    math_adder_full FA_13_04 (
        .i_a(w_sum_13_12),
        .i_b(w_sum_13_10),
        .i_c(w_sum_13_08),
        .ow_sum(w_sum_13_04),
        .ow_carry(w_carry_13_04)
    );
    wire w_sum_13_02, w_carry_13_02;
    math_adder_half HA_13_02 (
        .i_a(w_sum_13_06),
        .i_b(w_sum_13_04),
        .ow_sum(w_sum_13_02),
        .ow_carry(w_carry_13_02)
    );
    wire w_sum_14_28, w_carry_14_28;

    math_adder_full FA_14_28 (
        .i_a(w_pp_00_14),
        .i_b(w_pp_01_13),
        .i_c(w_pp_02_12),
        .ow_sum(w_sum_14_28),
        .ow_carry(w_carry_14_28)
    );
    wire w_sum_14_26, w_carry_14_26;

    math_adder_full FA_14_26 (
        .i_a(w_pp_03_11),
        .i_b(w_pp_04_10),
        .i_c(w_pp_05_09),
        .ow_sum(w_sum_14_26),
        .ow_carry(w_carry_14_26)
    );
    wire w_sum_14_24, w_carry_14_24;

    math_adder_full FA_14_24 (
        .i_a(w_pp_06_08),
        .i_b(w_pp_07_07),
        .i_c(w_pp_08_06),
        .ow_sum(w_sum_14_24),
        .ow_carry(w_carry_14_24)
    );
    wire w_sum_14_22, w_carry_14_22;

    math_adder_full FA_14_22 (
        .i_a(w_pp_09_05),
        .i_b(w_pp_10_04),
        .i_c(w_pp_11_03),
        .ow_sum(w_sum_14_22),
        .ow_carry(w_carry_14_22)
    );
    wire w_sum_14_20, w_carry_14_20;

    math_adder_full FA_14_20 (
        .i_a(w_pp_12_02),
        .i_b(w_pp_13_01),
        .i_c(w_pp_14_00),
        .ow_sum(w_sum_14_20),
        .ow_carry(w_carry_14_20)
    );
    wire w_sum_14_18, w_carry_14_18;

    math_adder_full FA_14_18 (
        .i_a(w_carry_13_26),
        .i_b(w_carry_13_24),
        .i_c(w_carry_13_22),
        .ow_sum(w_sum_14_18),
        .ow_carry(w_carry_14_18)
    );
    wire w_sum_14_16, w_carry_14_16;

    math_adder_full FA_14_16 (
        .i_a(w_carry_13_20),
        .i_b(w_carry_13_18),
        .i_c(w_carry_13_16),
        .ow_sum(w_sum_14_16),
        .ow_carry(w_carry_14_16)
    );
    wire w_sum_14_14, w_carry_14_14;

    math_adder_full FA_14_14 (
        .i_a(w_carry_13_14),
        .i_b(w_carry_13_12),
        .i_c(w_carry_13_10),
        .ow_sum(w_sum_14_14),
        .ow_carry(w_carry_14_14)
    );
    wire w_sum_14_12, w_carry_14_12;

    math_adder_full FA_14_12 (
        .i_a(w_carry_13_08),
        .i_b(w_carry_13_06),
        .i_c(w_carry_13_04),
        .ow_sum(w_sum_14_12),
        .ow_carry(w_carry_14_12)
    );
    wire w_sum_14_10, w_carry_14_10;

    math_adder_full FA_14_10 (
        .i_a(w_carry_13_02),
        .i_b(w_sum_14_28),
        .i_c(w_sum_14_26),
        .ow_sum(w_sum_14_10),
        .ow_carry(w_carry_14_10)
    );
    wire w_sum_14_08, w_carry_14_08;

    math_adder_full FA_14_08 (
        .i_a(w_sum_14_24),
        .i_b(w_sum_14_22),
        .i_c(w_sum_14_20),
        .ow_sum(w_sum_14_08),
        .ow_carry(w_carry_14_08)
    );
    wire w_sum_14_06, w_carry_14_06;

    math_adder_full FA_14_06 (
        .i_a(w_sum_14_18),
        .i_b(w_sum_14_16),
        .i_c(w_sum_14_14),
        .ow_sum(w_sum_14_06),
        .ow_carry(w_carry_14_06)
    );
    wire w_sum_14_04, w_carry_14_04;

    math_adder_full FA_14_04 (
        .i_a(w_sum_14_12),
        .i_b(w_sum_14_10),
        .i_c(w_sum_14_08),
        .ow_sum(w_sum_14_04),
        .ow_carry(w_carry_14_04)
    );
    wire w_sum_14_02, w_carry_14_02;
    math_adder_half HA_14_02 (
        .i_a(w_sum_14_06),
        .i_b(w_sum_14_04),
        .ow_sum(w_sum_14_02),
        .ow_carry(w_carry_14_02)
    );
    wire w_sum_15_30, w_carry_15_30;

    math_adder_full FA_15_30 (
        .i_a(w_pp_00_15),
        .i_b(w_pp_01_14),
        .i_c(w_pp_02_13),
        .ow_sum(w_sum_15_30),
        .ow_carry(w_carry_15_30)
    );
    wire w_sum_15_28, w_carry_15_28;

    math_adder_full FA_15_28 (
        .i_a(w_pp_03_12),
        .i_b(w_pp_04_11),
        .i_c(w_pp_05_10),
        .ow_sum(w_sum_15_28),
        .ow_carry(w_carry_15_28)
    );
    wire w_sum_15_26, w_carry_15_26;

    math_adder_full FA_15_26 (
        .i_a(w_pp_06_09),
        .i_b(w_pp_07_08),
        .i_c(w_pp_08_07),
        .ow_sum(w_sum_15_26),
        .ow_carry(w_carry_15_26)
    );
    wire w_sum_15_24, w_carry_15_24;

    math_adder_full FA_15_24 (
        .i_a(w_pp_09_06),
        .i_b(w_pp_10_05),
        .i_c(w_pp_11_04),
        .ow_sum(w_sum_15_24),
        .ow_carry(w_carry_15_24)
    );
    wire w_sum_15_22, w_carry_15_22;

    math_adder_full FA_15_22 (
        .i_a(w_pp_12_03),
        .i_b(w_pp_13_02),
        .i_c(w_pp_14_01),
        .ow_sum(w_sum_15_22),
        .ow_carry(w_carry_15_22)
    );
    wire w_sum_15_20, w_carry_15_20;

    math_adder_full FA_15_20 (
        .i_a(w_pp_15_00),
        .i_b(w_carry_14_28),
        .i_c(w_carry_14_26),
        .ow_sum(w_sum_15_20),
        .ow_carry(w_carry_15_20)
    );
    wire w_sum_15_18, w_carry_15_18;

    math_adder_full FA_15_18 (
        .i_a(w_carry_14_24),
        .i_b(w_carry_14_22),
        .i_c(w_carry_14_20),
        .ow_sum(w_sum_15_18),
        .ow_carry(w_carry_15_18)
    );
    wire w_sum_15_16, w_carry_15_16;

    math_adder_full FA_15_16 (
        .i_a(w_carry_14_18),
        .i_b(w_carry_14_16),
        .i_c(w_carry_14_14),
        .ow_sum(w_sum_15_16),
        .ow_carry(w_carry_15_16)
    );
    wire w_sum_15_14, w_carry_15_14;

    math_adder_full FA_15_14 (
        .i_a(w_carry_14_12),
        .i_b(w_carry_14_10),
        .i_c(w_carry_14_08),
        .ow_sum(w_sum_15_14),
        .ow_carry(w_carry_15_14)
    );
    wire w_sum_15_12, w_carry_15_12;

    math_adder_full FA_15_12 (
        .i_a(w_carry_14_06),
        .i_b(w_carry_14_04),
        .i_c(w_carry_14_02),
        .ow_sum(w_sum_15_12),
        .ow_carry(w_carry_15_12)
    );
    wire w_sum_15_10, w_carry_15_10;

    math_adder_full FA_15_10 (
        .i_a(w_sum_15_30),
        .i_b(w_sum_15_28),
        .i_c(w_sum_15_26),
        .ow_sum(w_sum_15_10),
        .ow_carry(w_carry_15_10)
    );
    wire w_sum_15_08, w_carry_15_08;

    math_adder_full FA_15_08 (
        .i_a(w_sum_15_24),
        .i_b(w_sum_15_22),
        .i_c(w_sum_15_20),
        .ow_sum(w_sum_15_08),
        .ow_carry(w_carry_15_08)
    );
    wire w_sum_15_06, w_carry_15_06;

    math_adder_full FA_15_06 (
        .i_a(w_sum_15_18),
        .i_b(w_sum_15_16),
        .i_c(w_sum_15_14),
        .ow_sum(w_sum_15_06),
        .ow_carry(w_carry_15_06)
    );
    wire w_sum_15_04, w_carry_15_04;

    math_adder_full FA_15_04 (
        .i_a(w_sum_15_12),
        .i_b(w_sum_15_10),
        .i_c(w_sum_15_08),
        .ow_sum(w_sum_15_04),
        .ow_carry(w_carry_15_04)
    );
    wire w_sum_15_02, w_carry_15_02;
    math_adder_half HA_15_02 (
        .i_a(w_sum_15_06),
        .i_b(w_sum_15_04),
        .ow_sum(w_sum_15_02),
        .ow_carry(w_carry_15_02)
    );
    wire w_sum_16_30, w_carry_16_30;

    math_adder_full FA_16_30 (
        .i_a(w_pp_01_15),
        .i_b(w_pp_02_14),
        .i_c(w_pp_03_13),
        .ow_sum(w_sum_16_30),
        .ow_carry(w_carry_16_30)
    );
    wire w_sum_16_28, w_carry_16_28;

    math_adder_full FA_16_28 (
        .i_a(w_pp_04_12),
        .i_b(w_pp_05_11),
        .i_c(w_pp_06_10),
        .ow_sum(w_sum_16_28),
        .ow_carry(w_carry_16_28)
    );
    wire w_sum_16_26, w_carry_16_26;

    math_adder_full FA_16_26 (
        .i_a(w_pp_07_09),
        .i_b(w_pp_08_08),
        .i_c(w_pp_09_07),
        .ow_sum(w_sum_16_26),
        .ow_carry(w_carry_16_26)
    );
    wire w_sum_16_24, w_carry_16_24;

    math_adder_full FA_16_24 (
        .i_a(w_pp_10_06),
        .i_b(w_pp_11_05),
        .i_c(w_pp_12_04),
        .ow_sum(w_sum_16_24),
        .ow_carry(w_carry_16_24)
    );
    wire w_sum_16_22, w_carry_16_22;

    math_adder_full FA_16_22 (
        .i_a(w_pp_13_03),
        .i_b(w_pp_14_02),
        .i_c(w_pp_15_01),
        .ow_sum(w_sum_16_22),
        .ow_carry(w_carry_16_22)
    );
    wire w_sum_16_20, w_carry_16_20;

    math_adder_full FA_16_20 (
        .i_a(w_carry_15_30),
        .i_b(w_carry_15_28),
        .i_c(w_carry_15_26),
        .ow_sum(w_sum_16_20),
        .ow_carry(w_carry_16_20)
    );
    wire w_sum_16_18, w_carry_16_18;

    math_adder_full FA_16_18 (
        .i_a(w_carry_15_24),
        .i_b(w_carry_15_22),
        .i_c(w_carry_15_20),
        .ow_sum(w_sum_16_18),
        .ow_carry(w_carry_16_18)
    );
    wire w_sum_16_16, w_carry_16_16;

    math_adder_full FA_16_16 (
        .i_a(w_carry_15_18),
        .i_b(w_carry_15_16),
        .i_c(w_carry_15_14),
        .ow_sum(w_sum_16_16),
        .ow_carry(w_carry_16_16)
    );
    wire w_sum_16_14, w_carry_16_14;

    math_adder_full FA_16_14 (
        .i_a(w_carry_15_12),
        .i_b(w_carry_15_10),
        .i_c(w_carry_15_08),
        .ow_sum(w_sum_16_14),
        .ow_carry(w_carry_16_14)
    );
    wire w_sum_16_12, w_carry_16_12;

    math_adder_full FA_16_12 (
        .i_a(w_carry_15_06),
        .i_b(w_carry_15_04),
        .i_c(w_carry_15_02),
        .ow_sum(w_sum_16_12),
        .ow_carry(w_carry_16_12)
    );
    wire w_sum_16_10, w_carry_16_10;

    math_adder_full FA_16_10 (
        .i_a(w_sum_16_30),
        .i_b(w_sum_16_28),
        .i_c(w_sum_16_26),
        .ow_sum(w_sum_16_10),
        .ow_carry(w_carry_16_10)
    );
    wire w_sum_16_08, w_carry_16_08;

    math_adder_full FA_16_08 (
        .i_a(w_sum_16_24),
        .i_b(w_sum_16_22),
        .i_c(w_sum_16_20),
        .ow_sum(w_sum_16_08),
        .ow_carry(w_carry_16_08)
    );
    wire w_sum_16_06, w_carry_16_06;

    math_adder_full FA_16_06 (
        .i_a(w_sum_16_18),
        .i_b(w_sum_16_16),
        .i_c(w_sum_16_14),
        .ow_sum(w_sum_16_06),
        .ow_carry(w_carry_16_06)
    );
    wire w_sum_16_04, w_carry_16_04;

    math_adder_full FA_16_04 (
        .i_a(w_sum_16_12),
        .i_b(w_sum_16_10),
        .i_c(w_sum_16_08),
        .ow_sum(w_sum_16_04),
        .ow_carry(w_carry_16_04)
    );
    wire w_sum_16_02, w_carry_16_02;
    math_adder_half HA_16_02 (
        .i_a(w_sum_16_06),
        .i_b(w_sum_16_04),
        .ow_sum(w_sum_16_02),
        .ow_carry(w_carry_16_02)
    );
    wire w_sum_17_29, w_carry_17_29;

    math_adder_full FA_17_29 (
        .i_a(w_pp_02_15),
        .i_b(w_pp_03_14),
        .i_c(w_pp_04_13),
        .ow_sum(w_sum_17_29),
        .ow_carry(w_carry_17_29)
    );
    wire w_sum_17_27, w_carry_17_27;

    math_adder_full FA_17_27 (
        .i_a(w_pp_05_12),
        .i_b(w_pp_06_11),
        .i_c(w_pp_07_10),
        .ow_sum(w_sum_17_27),
        .ow_carry(w_carry_17_27)
    );
    wire w_sum_17_25, w_carry_17_25;

    math_adder_full FA_17_25 (
        .i_a(w_pp_08_09),
        .i_b(w_pp_09_08),
        .i_c(w_pp_10_07),
        .ow_sum(w_sum_17_25),
        .ow_carry(w_carry_17_25)
    );
    wire w_sum_17_23, w_carry_17_23;

    math_adder_full FA_17_23 (
        .i_a(w_pp_11_06),
        .i_b(w_pp_12_05),
        .i_c(w_pp_13_04),
        .ow_sum(w_sum_17_23),
        .ow_carry(w_carry_17_23)
    );
    wire w_sum_17_21, w_carry_17_21;

    math_adder_full FA_17_21 (
        .i_a(w_pp_14_03),
        .i_b(w_pp_15_02),
        .i_c(w_carry_16_30),
        .ow_sum(w_sum_17_21),
        .ow_carry(w_carry_17_21)
    );
    wire w_sum_17_19, w_carry_17_19;

    math_adder_full FA_17_19 (
        .i_a(w_carry_16_28),
        .i_b(w_carry_16_26),
        .i_c(w_carry_16_24),
        .ow_sum(w_sum_17_19),
        .ow_carry(w_carry_17_19)
    );
    wire w_sum_17_17, w_carry_17_17;

    math_adder_full FA_17_17 (
        .i_a(w_carry_16_22),
        .i_b(w_carry_16_20),
        .i_c(w_carry_16_18),
        .ow_sum(w_sum_17_17),
        .ow_carry(w_carry_17_17)
    );
    wire w_sum_17_15, w_carry_17_15;

    math_adder_full FA_17_15 (
        .i_a(w_carry_16_16),
        .i_b(w_carry_16_14),
        .i_c(w_carry_16_12),
        .ow_sum(w_sum_17_15),
        .ow_carry(w_carry_17_15)
    );
    wire w_sum_17_13, w_carry_17_13;

    math_adder_full FA_17_13 (
        .i_a(w_carry_16_10),
        .i_b(w_carry_16_08),
        .i_c(w_carry_16_06),
        .ow_sum(w_sum_17_13),
        .ow_carry(w_carry_17_13)
    );
    wire w_sum_17_11, w_carry_17_11;

    math_adder_full FA_17_11 (
        .i_a(w_carry_16_04),
        .i_b(w_carry_16_02),
        .i_c(w_sum_17_29),
        .ow_sum(w_sum_17_11),
        .ow_carry(w_carry_17_11)
    );
    wire w_sum_17_09, w_carry_17_09;

    math_adder_full FA_17_09 (
        .i_a(w_sum_17_27),
        .i_b(w_sum_17_25),
        .i_c(w_sum_17_23),
        .ow_sum(w_sum_17_09),
        .ow_carry(w_carry_17_09)
    );
    wire w_sum_17_07, w_carry_17_07;

    math_adder_full FA_17_07 (
        .i_a(w_sum_17_21),
        .i_b(w_sum_17_19),
        .i_c(w_sum_17_17),
        .ow_sum(w_sum_17_07),
        .ow_carry(w_carry_17_07)
    );
    wire w_sum_17_05, w_carry_17_05;

    math_adder_full FA_17_05 (
        .i_a(w_sum_17_15),
        .i_b(w_sum_17_13),
        .i_c(w_sum_17_11),
        .ow_sum(w_sum_17_05),
        .ow_carry(w_carry_17_05)
    );
    wire w_sum_17_03, w_carry_17_03;

    math_adder_full FA_17_03 (
        .i_a(w_sum_17_09),
        .i_b(w_sum_17_07),
        .i_c(w_sum_17_05),
        .ow_sum(w_sum_17_03),
        .ow_carry(w_carry_17_03)
    );
    wire w_sum_18_27, w_carry_18_27;

    math_adder_full FA_18_27 (
        .i_a(w_pp_03_15),
        .i_b(w_pp_04_14),
        .i_c(w_pp_05_13),
        .ow_sum(w_sum_18_27),
        .ow_carry(w_carry_18_27)
    );
    wire w_sum_18_25, w_carry_18_25;

    math_adder_full FA_18_25 (
        .i_a(w_pp_06_12),
        .i_b(w_pp_07_11),
        .i_c(w_pp_08_10),
        .ow_sum(w_sum_18_25),
        .ow_carry(w_carry_18_25)
    );
    wire w_sum_18_23, w_carry_18_23;

    math_adder_full FA_18_23 (
        .i_a(w_pp_09_09),
        .i_b(w_pp_10_08),
        .i_c(w_pp_11_07),
        .ow_sum(w_sum_18_23),
        .ow_carry(w_carry_18_23)
    );
    wire w_sum_18_21, w_carry_18_21;

    math_adder_full FA_18_21 (
        .i_a(w_pp_12_06),
        .i_b(w_pp_13_05),
        .i_c(w_pp_14_04),
        .ow_sum(w_sum_18_21),
        .ow_carry(w_carry_18_21)
    );
    wire w_sum_18_19, w_carry_18_19;

    math_adder_full FA_18_19 (
        .i_a(w_pp_15_03),
        .i_b(w_carry_17_29),
        .i_c(w_carry_17_27),
        .ow_sum(w_sum_18_19),
        .ow_carry(w_carry_18_19)
    );
    wire w_sum_18_17, w_carry_18_17;

    math_adder_full FA_18_17 (
        .i_a(w_carry_17_25),
        .i_b(w_carry_17_23),
        .i_c(w_carry_17_21),
        .ow_sum(w_sum_18_17),
        .ow_carry(w_carry_18_17)
    );
    wire w_sum_18_15, w_carry_18_15;

    math_adder_full FA_18_15 (
        .i_a(w_carry_17_19),
        .i_b(w_carry_17_17),
        .i_c(w_carry_17_15),
        .ow_sum(w_sum_18_15),
        .ow_carry(w_carry_18_15)
    );
    wire w_sum_18_13, w_carry_18_13;

    math_adder_full FA_18_13 (
        .i_a(w_carry_17_13),
        .i_b(w_carry_17_11),
        .i_c(w_carry_17_09),
        .ow_sum(w_sum_18_13),
        .ow_carry(w_carry_18_13)
    );
    wire w_sum_18_11, w_carry_18_11;

    math_adder_full FA_18_11 (
        .i_a(w_carry_17_07),
        .i_b(w_carry_17_05),
        .i_c(w_carry_17_03),
        .ow_sum(w_sum_18_11),
        .ow_carry(w_carry_18_11)
    );
    wire w_sum_18_09, w_carry_18_09;

    math_adder_full FA_18_09 (
        .i_a(w_sum_18_27),
        .i_b(w_sum_18_25),
        .i_c(w_sum_18_23),
        .ow_sum(w_sum_18_09),
        .ow_carry(w_carry_18_09)
    );
    wire w_sum_18_07, w_carry_18_07;

    math_adder_full FA_18_07 (
        .i_a(w_sum_18_21),
        .i_b(w_sum_18_19),
        .i_c(w_sum_18_17),
        .ow_sum(w_sum_18_07),
        .ow_carry(w_carry_18_07)
    );
    wire w_sum_18_05, w_carry_18_05;

    math_adder_full FA_18_05 (
        .i_a(w_sum_18_15),
        .i_b(w_sum_18_13),
        .i_c(w_sum_18_11),
        .ow_sum(w_sum_18_05),
        .ow_carry(w_carry_18_05)
    );
    wire w_sum_18_03, w_carry_18_03;

    math_adder_full FA_18_03 (
        .i_a(w_sum_18_09),
        .i_b(w_sum_18_07),
        .i_c(w_sum_18_05),
        .ow_sum(w_sum_18_03),
        .ow_carry(w_carry_18_03)
    );
    wire w_sum_19_25, w_carry_19_25;

    math_adder_full FA_19_25 (
        .i_a(w_pp_04_15),
        .i_b(w_pp_05_14),
        .i_c(w_pp_06_13),
        .ow_sum(w_sum_19_25),
        .ow_carry(w_carry_19_25)
    );
    wire w_sum_19_23, w_carry_19_23;

    math_adder_full FA_19_23 (
        .i_a(w_pp_07_12),
        .i_b(w_pp_08_11),
        .i_c(w_pp_09_10),
        .ow_sum(w_sum_19_23),
        .ow_carry(w_carry_19_23)
    );
    wire w_sum_19_21, w_carry_19_21;

    math_adder_full FA_19_21 (
        .i_a(w_pp_10_09),
        .i_b(w_pp_11_08),
        .i_c(w_pp_12_07),
        .ow_sum(w_sum_19_21),
        .ow_carry(w_carry_19_21)
    );
    wire w_sum_19_19, w_carry_19_19;

    math_adder_full FA_19_19 (
        .i_a(w_pp_13_06),
        .i_b(w_pp_14_05),
        .i_c(w_pp_15_04),
        .ow_sum(w_sum_19_19),
        .ow_carry(w_carry_19_19)
    );
    wire w_sum_19_17, w_carry_19_17;

    math_adder_full FA_19_17 (
        .i_a(w_carry_18_27),
        .i_b(w_carry_18_25),
        .i_c(w_carry_18_23),
        .ow_sum(w_sum_19_17),
        .ow_carry(w_carry_19_17)
    );
    wire w_sum_19_15, w_carry_19_15;

    math_adder_full FA_19_15 (
        .i_a(w_carry_18_21),
        .i_b(w_carry_18_19),
        .i_c(w_carry_18_17),
        .ow_sum(w_sum_19_15),
        .ow_carry(w_carry_19_15)
    );
    wire w_sum_19_13, w_carry_19_13;

    math_adder_full FA_19_13 (
        .i_a(w_carry_18_15),
        .i_b(w_carry_18_13),
        .i_c(w_carry_18_11),
        .ow_sum(w_sum_19_13),
        .ow_carry(w_carry_19_13)
    );
    wire w_sum_19_11, w_carry_19_11;

    math_adder_full FA_19_11 (
        .i_a(w_carry_18_09),
        .i_b(w_carry_18_07),
        .i_c(w_carry_18_05),
        .ow_sum(w_sum_19_11),
        .ow_carry(w_carry_19_11)
    );
    wire w_sum_19_09, w_carry_19_09;

    math_adder_full FA_19_09 (
        .i_a(w_carry_18_03),
        .i_b(w_sum_19_25),
        .i_c(w_sum_19_23),
        .ow_sum(w_sum_19_09),
        .ow_carry(w_carry_19_09)
    );
    wire w_sum_19_07, w_carry_19_07;

    math_adder_full FA_19_07 (
        .i_a(w_sum_19_21),
        .i_b(w_sum_19_19),
        .i_c(w_sum_19_17),
        .ow_sum(w_sum_19_07),
        .ow_carry(w_carry_19_07)
    );
    wire w_sum_19_05, w_carry_19_05;

    math_adder_full FA_19_05 (
        .i_a(w_sum_19_15),
        .i_b(w_sum_19_13),
        .i_c(w_sum_19_11),
        .ow_sum(w_sum_19_05),
        .ow_carry(w_carry_19_05)
    );
    wire w_sum_19_03, w_carry_19_03;

    math_adder_full FA_19_03 (
        .i_a(w_sum_19_09),
        .i_b(w_sum_19_07),
        .i_c(w_sum_19_05),
        .ow_sum(w_sum_19_03),
        .ow_carry(w_carry_19_03)
    );
    wire w_sum_20_23, w_carry_20_23;

    math_adder_full FA_20_23 (
        .i_a(w_pp_05_15),
        .i_b(w_pp_06_14),
        .i_c(w_pp_07_13),
        .ow_sum(w_sum_20_23),
        .ow_carry(w_carry_20_23)
    );
    wire w_sum_20_21, w_carry_20_21;

    math_adder_full FA_20_21 (
        .i_a(w_pp_08_12),
        .i_b(w_pp_09_11),
        .i_c(w_pp_10_10),
        .ow_sum(w_sum_20_21),
        .ow_carry(w_carry_20_21)
    );
    wire w_sum_20_19, w_carry_20_19;

    math_adder_full FA_20_19 (
        .i_a(w_pp_11_09),
        .i_b(w_pp_12_08),
        .i_c(w_pp_13_07),
        .ow_sum(w_sum_20_19),
        .ow_carry(w_carry_20_19)
    );
    wire w_sum_20_17, w_carry_20_17;

    math_adder_full FA_20_17 (
        .i_a(w_pp_14_06),
        .i_b(w_pp_15_05),
        .i_c(w_carry_19_25),
        .ow_sum(w_sum_20_17),
        .ow_carry(w_carry_20_17)
    );
    wire w_sum_20_15, w_carry_20_15;

    math_adder_full FA_20_15 (
        .i_a(w_carry_19_23),
        .i_b(w_carry_19_21),
        .i_c(w_carry_19_19),
        .ow_sum(w_sum_20_15),
        .ow_carry(w_carry_20_15)
    );
    wire w_sum_20_13, w_carry_20_13;

    math_adder_full FA_20_13 (
        .i_a(w_carry_19_17),
        .i_b(w_carry_19_15),
        .i_c(w_carry_19_13),
        .ow_sum(w_sum_20_13),
        .ow_carry(w_carry_20_13)
    );
    wire w_sum_20_11, w_carry_20_11;

    math_adder_full FA_20_11 (
        .i_a(w_carry_19_11),
        .i_b(w_carry_19_09),
        .i_c(w_carry_19_07),
        .ow_sum(w_sum_20_11),
        .ow_carry(w_carry_20_11)
    );
    wire w_sum_20_09, w_carry_20_09;

    math_adder_full FA_20_09 (
        .i_a(w_carry_19_05),
        .i_b(w_carry_19_03),
        .i_c(w_sum_20_23),
        .ow_sum(w_sum_20_09),
        .ow_carry(w_carry_20_09)
    );
    wire w_sum_20_07, w_carry_20_07;

    math_adder_full FA_20_07 (
        .i_a(w_sum_20_21),
        .i_b(w_sum_20_19),
        .i_c(w_sum_20_17),
        .ow_sum(w_sum_20_07),
        .ow_carry(w_carry_20_07)
    );
    wire w_sum_20_05, w_carry_20_05;

    math_adder_full FA_20_05 (
        .i_a(w_sum_20_15),
        .i_b(w_sum_20_13),
        .i_c(w_sum_20_11),
        .ow_sum(w_sum_20_05),
        .ow_carry(w_carry_20_05)
    );
    wire w_sum_20_03, w_carry_20_03;

    math_adder_full FA_20_03 (
        .i_a(w_sum_20_09),
        .i_b(w_sum_20_07),
        .i_c(w_sum_20_05),
        .ow_sum(w_sum_20_03),
        .ow_carry(w_carry_20_03)
    );
    wire w_sum_21_21, w_carry_21_21;

    math_adder_full FA_21_21 (
        .i_a(w_pp_06_15),
        .i_b(w_pp_07_14),
        .i_c(w_pp_08_13),
        .ow_sum(w_sum_21_21),
        .ow_carry(w_carry_21_21)
    );
    wire w_sum_21_19, w_carry_21_19;

    math_adder_full FA_21_19 (
        .i_a(w_pp_09_12),
        .i_b(w_pp_10_11),
        .i_c(w_pp_11_10),
        .ow_sum(w_sum_21_19),
        .ow_carry(w_carry_21_19)
    );
    wire w_sum_21_17, w_carry_21_17;

    math_adder_full FA_21_17 (
        .i_a(w_pp_12_09),
        .i_b(w_pp_13_08),
        .i_c(w_pp_14_07),
        .ow_sum(w_sum_21_17),
        .ow_carry(w_carry_21_17)
    );
    wire w_sum_21_15, w_carry_21_15;

    math_adder_full FA_21_15 (
        .i_a(w_pp_15_06),
        .i_b(w_carry_20_23),
        .i_c(w_carry_20_21),
        .ow_sum(w_sum_21_15),
        .ow_carry(w_carry_21_15)
    );
    wire w_sum_21_13, w_carry_21_13;

    math_adder_full FA_21_13 (
        .i_a(w_carry_20_19),
        .i_b(w_carry_20_17),
        .i_c(w_carry_20_15),
        .ow_sum(w_sum_21_13),
        .ow_carry(w_carry_21_13)
    );
    wire w_sum_21_11, w_carry_21_11;

    math_adder_full FA_21_11 (
        .i_a(w_carry_20_13),
        .i_b(w_carry_20_11),
        .i_c(w_carry_20_09),
        .ow_sum(w_sum_21_11),
        .ow_carry(w_carry_21_11)
    );
    wire w_sum_21_09, w_carry_21_09;

    math_adder_full FA_21_09 (
        .i_a(w_carry_20_07),
        .i_b(w_carry_20_05),
        .i_c(w_carry_20_03),
        .ow_sum(w_sum_21_09),
        .ow_carry(w_carry_21_09)
    );
    wire w_sum_21_07, w_carry_21_07;

    math_adder_full FA_21_07 (
        .i_a(w_sum_21_21),
        .i_b(w_sum_21_19),
        .i_c(w_sum_21_17),
        .ow_sum(w_sum_21_07),
        .ow_carry(w_carry_21_07)
    );
    wire w_sum_21_05, w_carry_21_05;

    math_adder_full FA_21_05 (
        .i_a(w_sum_21_15),
        .i_b(w_sum_21_13),
        .i_c(w_sum_21_11),
        .ow_sum(w_sum_21_05),
        .ow_carry(w_carry_21_05)
    );
    wire w_sum_21_03, w_carry_21_03;

    math_adder_full FA_21_03 (
        .i_a(w_sum_21_09),
        .i_b(w_sum_21_07),
        .i_c(w_sum_21_05),
        .ow_sum(w_sum_21_03),
        .ow_carry(w_carry_21_03)
    );
    wire w_sum_22_19, w_carry_22_19;

    math_adder_full FA_22_19 (
        .i_a(w_pp_07_15),
        .i_b(w_pp_08_14),
        .i_c(w_pp_09_13),
        .ow_sum(w_sum_22_19),
        .ow_carry(w_carry_22_19)
    );
    wire w_sum_22_17, w_carry_22_17;

    math_adder_full FA_22_17 (
        .i_a(w_pp_10_12),
        .i_b(w_pp_11_11),
        .i_c(w_pp_12_10),
        .ow_sum(w_sum_22_17),
        .ow_carry(w_carry_22_17)
    );
    wire w_sum_22_15, w_carry_22_15;

    math_adder_full FA_22_15 (
        .i_a(w_pp_13_09),
        .i_b(w_pp_14_08),
        .i_c(w_pp_15_07),
        .ow_sum(w_sum_22_15),
        .ow_carry(w_carry_22_15)
    );
    wire w_sum_22_13, w_carry_22_13;

    math_adder_full FA_22_13 (
        .i_a(w_carry_21_21),
        .i_b(w_carry_21_19),
        .i_c(w_carry_21_17),
        .ow_sum(w_sum_22_13),
        .ow_carry(w_carry_22_13)
    );
    wire w_sum_22_11, w_carry_22_11;

    math_adder_full FA_22_11 (
        .i_a(w_carry_21_15),
        .i_b(w_carry_21_13),
        .i_c(w_carry_21_11),
        .ow_sum(w_sum_22_11),
        .ow_carry(w_carry_22_11)
    );
    wire w_sum_22_09, w_carry_22_09;

    math_adder_full FA_22_09 (
        .i_a(w_carry_21_09),
        .i_b(w_carry_21_07),
        .i_c(w_carry_21_05),
        .ow_sum(w_sum_22_09),
        .ow_carry(w_carry_22_09)
    );
    wire w_sum_22_07, w_carry_22_07;

    math_adder_full FA_22_07 (
        .i_a(w_carry_21_03),
        .i_b(w_sum_22_19),
        .i_c(w_sum_22_17),
        .ow_sum(w_sum_22_07),
        .ow_carry(w_carry_22_07)
    );
    wire w_sum_22_05, w_carry_22_05;

    math_adder_full FA_22_05 (
        .i_a(w_sum_22_15),
        .i_b(w_sum_22_13),
        .i_c(w_sum_22_11),
        .ow_sum(w_sum_22_05),
        .ow_carry(w_carry_22_05)
    );
    wire w_sum_22_03, w_carry_22_03;

    math_adder_full FA_22_03 (
        .i_a(w_sum_22_09),
        .i_b(w_sum_22_07),
        .i_c(w_sum_22_05),
        .ow_sum(w_sum_22_03),
        .ow_carry(w_carry_22_03)
    );
    wire w_sum_23_17, w_carry_23_17;

    math_adder_full FA_23_17 (
        .i_a(w_pp_08_15),
        .i_b(w_pp_09_14),
        .i_c(w_pp_10_13),
        .ow_sum(w_sum_23_17),
        .ow_carry(w_carry_23_17)
    );
    wire w_sum_23_15, w_carry_23_15;

    math_adder_full FA_23_15 (
        .i_a(w_pp_11_12),
        .i_b(w_pp_12_11),
        .i_c(w_pp_13_10),
        .ow_sum(w_sum_23_15),
        .ow_carry(w_carry_23_15)
    );
    wire w_sum_23_13, w_carry_23_13;

    math_adder_full FA_23_13 (
        .i_a(w_pp_14_09),
        .i_b(w_pp_15_08),
        .i_c(w_carry_22_19),
        .ow_sum(w_sum_23_13),
        .ow_carry(w_carry_23_13)
    );
    wire w_sum_23_11, w_carry_23_11;

    math_adder_full FA_23_11 (
        .i_a(w_carry_22_17),
        .i_b(w_carry_22_15),
        .i_c(w_carry_22_13),
        .ow_sum(w_sum_23_11),
        .ow_carry(w_carry_23_11)
    );
    wire w_sum_23_09, w_carry_23_09;

    math_adder_full FA_23_09 (
        .i_a(w_carry_22_11),
        .i_b(w_carry_22_09),
        .i_c(w_carry_22_07),
        .ow_sum(w_sum_23_09),
        .ow_carry(w_carry_23_09)
    );
    wire w_sum_23_07, w_carry_23_07;

    math_adder_full FA_23_07 (
        .i_a(w_carry_22_05),
        .i_b(w_carry_22_03),
        .i_c(w_sum_23_17),
        .ow_sum(w_sum_23_07),
        .ow_carry(w_carry_23_07)
    );
    wire w_sum_23_05, w_carry_23_05;

    math_adder_full FA_23_05 (
        .i_a(w_sum_23_15),
        .i_b(w_sum_23_13),
        .i_c(w_sum_23_11),
        .ow_sum(w_sum_23_05),
        .ow_carry(w_carry_23_05)
    );
    wire w_sum_23_03, w_carry_23_03;

    math_adder_full FA_23_03 (
        .i_a(w_sum_23_09),
        .i_b(w_sum_23_07),
        .i_c(w_sum_23_05),
        .ow_sum(w_sum_23_03),
        .ow_carry(w_carry_23_03)
    );
    wire w_sum_24_15, w_carry_24_15;

    math_adder_full FA_24_15 (
        .i_a(w_pp_09_15),
        .i_b(w_pp_10_14),
        .i_c(w_pp_11_13),
        .ow_sum(w_sum_24_15),
        .ow_carry(w_carry_24_15)
    );
    wire w_sum_24_13, w_carry_24_13;

    math_adder_full FA_24_13 (
        .i_a(w_pp_12_12),
        .i_b(w_pp_13_11),
        .i_c(w_pp_14_10),
        .ow_sum(w_sum_24_13),
        .ow_carry(w_carry_24_13)
    );
    wire w_sum_24_11, w_carry_24_11;

    math_adder_full FA_24_11 (
        .i_a(w_pp_15_09),
        .i_b(w_carry_23_17),
        .i_c(w_carry_23_15),
        .ow_sum(w_sum_24_11),
        .ow_carry(w_carry_24_11)
    );
    wire w_sum_24_09, w_carry_24_09;

    math_adder_full FA_24_09 (
        .i_a(w_carry_23_13),
        .i_b(w_carry_23_11),
        .i_c(w_carry_23_09),
        .ow_sum(w_sum_24_09),
        .ow_carry(w_carry_24_09)
    );
    wire w_sum_24_07, w_carry_24_07;

    math_adder_full FA_24_07 (
        .i_a(w_carry_23_07),
        .i_b(w_carry_23_05),
        .i_c(w_carry_23_03),
        .ow_sum(w_sum_24_07),
        .ow_carry(w_carry_24_07)
    );
    wire w_sum_24_05, w_carry_24_05;

    math_adder_full FA_24_05 (
        .i_a(w_sum_24_15),
        .i_b(w_sum_24_13),
        .i_c(w_sum_24_11),
        .ow_sum(w_sum_24_05),
        .ow_carry(w_carry_24_05)
    );
    wire w_sum_24_03, w_carry_24_03;

    math_adder_full FA_24_03 (
        .i_a(w_sum_24_09),
        .i_b(w_sum_24_07),
        .i_c(w_sum_24_05),
        .ow_sum(w_sum_24_03),
        .ow_carry(w_carry_24_03)
    );
    wire w_sum_25_13, w_carry_25_13;

    math_adder_full FA_25_13 (
        .i_a(w_pp_10_15),
        .i_b(w_pp_11_14),
        .i_c(w_pp_12_13),
        .ow_sum(w_sum_25_13),
        .ow_carry(w_carry_25_13)
    );
    wire w_sum_25_11, w_carry_25_11;

    math_adder_full FA_25_11 (
        .i_a(w_pp_13_12),
        .i_b(w_pp_14_11),
        .i_c(w_pp_15_10),
        .ow_sum(w_sum_25_11),
        .ow_carry(w_carry_25_11)
    );
    wire w_sum_25_09, w_carry_25_09;

    math_adder_full FA_25_09 (
        .i_a(w_carry_24_15),
        .i_b(w_carry_24_13),
        .i_c(w_carry_24_11),
        .ow_sum(w_sum_25_09),
        .ow_carry(w_carry_25_09)
    );
    wire w_sum_25_07, w_carry_25_07;

    math_adder_full FA_25_07 (
        .i_a(w_carry_24_09),
        .i_b(w_carry_24_07),
        .i_c(w_carry_24_05),
        .ow_sum(w_sum_25_07),
        .ow_carry(w_carry_25_07)
    );
    wire w_sum_25_05, w_carry_25_05;

    math_adder_full FA_25_05 (
        .i_a(w_carry_24_03),
        .i_b(w_sum_25_13),
        .i_c(w_sum_25_11),
        .ow_sum(w_sum_25_05),
        .ow_carry(w_carry_25_05)
    );
    wire w_sum_25_03, w_carry_25_03;

    math_adder_full FA_25_03 (
        .i_a(w_sum_25_09),
        .i_b(w_sum_25_07),
        .i_c(w_sum_25_05),
        .ow_sum(w_sum_25_03),
        .ow_carry(w_carry_25_03)
    );
    wire w_sum_26_11, w_carry_26_11;

    math_adder_full FA_26_11 (
        .i_a(w_pp_11_15),
        .i_b(w_pp_12_14),
        .i_c(w_pp_13_13),
        .ow_sum(w_sum_26_11),
        .ow_carry(w_carry_26_11)
    );
    wire w_sum_26_09, w_carry_26_09;

    math_adder_full FA_26_09 (
        .i_a(w_pp_14_12),
        .i_b(w_pp_15_11),
        .i_c(w_carry_25_13),
        .ow_sum(w_sum_26_09),
        .ow_carry(w_carry_26_09)
    );
    wire w_sum_26_07, w_carry_26_07;

    math_adder_full FA_26_07 (
        .i_a(w_carry_25_11),
        .i_b(w_carry_25_09),
        .i_c(w_carry_25_07),
        .ow_sum(w_sum_26_07),
        .ow_carry(w_carry_26_07)
    );
    wire w_sum_26_05, w_carry_26_05;

    math_adder_full FA_26_05 (
        .i_a(w_carry_25_05),
        .i_b(w_carry_25_03),
        .i_c(w_sum_26_11),
        .ow_sum(w_sum_26_05),
        .ow_carry(w_carry_26_05)
    );
    wire w_sum_26_03, w_carry_26_03;

    math_adder_full FA_26_03 (
        .i_a(w_sum_26_09),
        .i_b(w_sum_26_07),
        .i_c(w_sum_26_05),
        .ow_sum(w_sum_26_03),
        .ow_carry(w_carry_26_03)
    );
    wire w_sum_27_09, w_carry_27_09;

    math_adder_full FA_27_09 (
        .i_a(w_pp_12_15),
        .i_b(w_pp_13_14),
        .i_c(w_pp_14_13),
        .ow_sum(w_sum_27_09),
        .ow_carry(w_carry_27_09)
    );
    wire w_sum_27_07, w_carry_27_07;

    math_adder_full FA_27_07 (
        .i_a(w_pp_15_12),
        .i_b(w_carry_26_11),
        .i_c(w_carry_26_09),
        .ow_sum(w_sum_27_07),
        .ow_carry(w_carry_27_07)
    );
    wire w_sum_27_05, w_carry_27_05;

    math_adder_full FA_27_05 (
        .i_a(w_carry_26_07),
        .i_b(w_carry_26_05),
        .i_c(w_carry_26_03),
        .ow_sum(w_sum_27_05),
        .ow_carry(w_carry_27_05)
    );
    wire w_sum_27_03, w_carry_27_03;

    math_adder_full FA_27_03 (
        .i_a(w_sum_27_09),
        .i_b(w_sum_27_07),
        .i_c(w_sum_27_05),
        .ow_sum(w_sum_27_03),
        .ow_carry(w_carry_27_03)
    );
    wire w_sum_28_07, w_carry_28_07;

    math_adder_full FA_28_07 (
        .i_a(w_pp_13_15),
        .i_b(w_pp_14_14),
        .i_c(w_pp_15_13),
        .ow_sum(w_sum_28_07),
        .ow_carry(w_carry_28_07)
    );
    wire w_sum_28_05, w_carry_28_05;

    math_adder_full FA_28_05 (
        .i_a(w_carry_27_09),
        .i_b(w_carry_27_07),
        .i_c(w_carry_27_05),
        .ow_sum(w_sum_28_05),
        .ow_carry(w_carry_28_05)
    );
    wire w_sum_28_03, w_carry_28_03;

    math_adder_full FA_28_03 (
        .i_a(w_carry_27_03),
        .i_b(w_sum_28_07),
        .i_c(w_sum_28_05),
        .ow_sum(w_sum_28_03),
        .ow_carry(w_carry_28_03)
    );
    wire w_sum_29_05, w_carry_29_05;

    math_adder_full FA_29_05 (
        .i_a(w_pp_14_15),
        .i_b(w_pp_15_14),
        .i_c(w_carry_28_07),
        .ow_sum(w_sum_29_05),
        .ow_carry(w_carry_29_05)
    );
    wire w_sum_29_03, w_carry_29_03;

    math_adder_full FA_29_03 (
        .i_a(w_carry_28_05),
        .i_b(w_carry_28_03),
        .i_c(w_sum_29_05),
        .ow_sum(w_sum_29_03),
        .ow_carry(w_carry_29_03)
    );
    wire w_sum_30_03, w_carry_30_03;

    math_adder_full FA_30_03 (
        .i_a(w_pp_15_15),
        .i_b(w_carry_29_05),
        .i_c(w_carry_29_03),
        .ow_sum(w_sum_30_03),
        .ow_carry(w_carry_30_03)
    );

    // Final addition stage
    wire w_sum_00 = w_pp_00_00;
    wire w_carry_00 = 1'b0;
    wire w_sum_01 = w_sum_01_02;
    wire w_carry_01 = 1'b0;
    wire w_sum_02 = w_sum_02_02;
    wire w_carry_02 = 1'b0;
    wire w_sum_03 = w_sum_03_02;
    wire w_carry_03 = 1'b0;
    wire w_sum_04 = w_sum_04_02;
    wire w_carry_04 = 1'b0;
    wire w_sum_05 = w_sum_05_02;
    wire w_carry_05 = 1'b0;
    wire w_sum_06 = w_sum_06_02;
    wire w_carry_06 = 1'b0;
    wire w_sum_07 = w_sum_07_02;
    wire w_carry_07 = 1'b0;
    wire w_sum_08 = w_sum_08_02;
    wire w_carry_08 = 1'b0;
    wire w_sum_09 = w_sum_09_02;
    wire w_carry_09 = 1'b0;
    wire w_sum_10 = w_sum_10_02;
    wire w_carry_10 = 1'b0;
    wire w_sum_11 = w_sum_11_02;
    wire w_carry_11 = 1'b0;
    wire w_sum_12 = w_sum_12_02;
    wire w_carry_12 = 1'b0;
    wire w_sum_13 = w_sum_13_02;
    wire w_carry_13 = 1'b0;
    wire w_sum_14 = w_sum_14_02;
    wire w_carry_14 = 1'b0;
    wire w_sum_15 = w_sum_15_02;
    wire w_carry_15 = 1'b0;
    wire w_sum_16 = w_sum_16_02;
    wire w_carry_16 = 1'b0;
    wire w_sum_17 = w_sum_17_03;
    wire w_carry_17 = 1'b0;
    wire w_sum_18 = w_sum_18_03;
    wire w_carry_18 = 1'b0;
    wire w_sum_19 = w_sum_19_03;
    wire w_carry_19 = 1'b0;
    wire w_sum_20 = w_sum_20_03;
    wire w_carry_20 = 1'b0;
    wire w_sum_21 = w_sum_21_03;
    wire w_carry_21 = 1'b0;
    wire w_sum_22 = w_sum_22_03;
    wire w_carry_22 = 1'b0;
    wire w_sum_23 = w_sum_23_03;
    wire w_carry_23 = 1'b0;
    wire w_sum_24 = w_sum_24_03;
    wire w_carry_24 = 1'b0;
    wire w_sum_25 = w_sum_25_03;
    wire w_carry_25 = 1'b0;
    wire w_sum_26 = w_sum_26_03;
    wire w_carry_26 = 1'b0;
    wire w_sum_27 = w_sum_27_03;
    wire w_carry_27 = 1'b0;
    wire w_sum_28 = w_sum_28_03;
    wire w_carry_28 = 1'b0;
    wire w_sum_29 = w_sum_29_03;
    wire w_carry_29 = 1'b0;
    wire w_sum_30 = w_sum_30_03;
    wire w_carry_30 = 1'b0;
    wire w_sum_31 = w_carry_30_03;
    wire w_carry_31 = 1'b0;

    // Final product assignment
    assign ow_product[0]  = w_sum_00;
    assign ow_product[1]  = w_sum_01;
    assign ow_product[2]  = w_sum_02;
    assign ow_product[3]  = w_sum_03;
    assign ow_product[4]  = w_sum_04;
    assign ow_product[5]  = w_sum_05;
    assign ow_product[6]  = w_sum_06;
    assign ow_product[7]  = w_sum_07;
    assign ow_product[8]  = w_sum_08;
    assign ow_product[9]  = w_sum_09;
    assign ow_product[10] = w_sum_10;
    assign ow_product[11] = w_sum_11;
    assign ow_product[12] = w_sum_12;
    assign ow_product[13] = w_sum_13;
    assign ow_product[14] = w_sum_14;
    assign ow_product[15] = w_sum_15;
    assign ow_product[16] = w_sum_16;
    assign ow_product[17] = w_sum_17;
    assign ow_product[18] = w_sum_18;
    assign ow_product[19] = w_sum_19;
    assign ow_product[20] = w_sum_20;
    assign ow_product[21] = w_sum_21;
    assign ow_product[22] = w_sum_22;
    assign ow_product[23] = w_sum_23;
    assign ow_product[24] = w_sum_24;
    assign ow_product[25] = w_sum_25;
    assign ow_product[26] = w_sum_26;
    assign ow_product[27] = w_sum_27;
    assign ow_product[28] = w_sum_28;
    assign ow_product[29] = w_sum_29;
    assign ow_product[30] = w_sum_30;
    assign ow_product[31] = w_sum_31;


    // synopsys translate_off
    initial begin
        $dumpfile("waves.vcd");
        $dumpvars(0, math_multiplier_wallace_tree_016);
    end
    // synopsys translate_on

endmodule
