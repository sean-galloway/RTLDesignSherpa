// SPDX-License-Identifier: MIT
// SPDX-FileCopyrightText: 2024-2025 sean galloway
//
// RTL Design Sherpa - Industry-Standard RTL Design and Verification
// https://github.com/sean-galloway/RTLDesignSherpa
//
// Module: bus_types
// Purpose: Bus Types module
//
// Documentation: rtl/amba/PRD.md
// Subsystem: amba
//
// Author: sean galloway
// Created: 2025-10-18

`ifndef BUS_TYPES_SVH
`define BUS_TYPES_SVH

`include "axi_pkg.sv"
`include "apb_pkg.sv"

`endif // BUS_TYPES_SVH
