// SPDX-License-Identifier: MIT
// SPDX-FileCopyrightText: 2024-2025 sean galloway
//
// RTL Design Sherpa - Industry-Standard RTL Design and Verification
// https://github.com/sean-galloway/RTLDesignSherpa
//
// Module: math_multiplier_dadda_4to2_024
// Purpose: Dadda 24x24 multiplier with 4:2 compressors for FP32 mantissa
//
// Documentation: IEEE754_ARCHITECTURE.md
// Subsystem: common
//
// Author: sean galloway
// Created: 2026-01-03
//
// AUTO-GENERATED FILE - DO NOT EDIT MANUALLY
// Generator: bin/rtl_generators/ieee754/dadda_4to2_multiplier.py
// Regenerate: PYTHONPATH=bin:$PYTHONPATH python3 bin/rtl_generators/ieee754/generate_all.py rtl/common
//

`timescale 1ns / 1ps

module math_multiplier_dadda_4to2_024 #(parameter int  N = 24)(
    input  logic [N-1:0]   i_multiplier,
    input  logic [N-1:0]   i_multiplicand,
    output logic [2*N-1:0] ow_product
);

// Partial Products (AND gate array)
wire w_pp_00_00 = i_multiplier[0] & i_multiplicand[0];
wire w_pp_00_01 = i_multiplier[0] & i_multiplicand[1];
wire w_pp_00_02 = i_multiplier[0] & i_multiplicand[2];
wire w_pp_00_03 = i_multiplier[0] & i_multiplicand[3];
wire w_pp_00_04 = i_multiplier[0] & i_multiplicand[4];
wire w_pp_00_05 = i_multiplier[0] & i_multiplicand[5];
wire w_pp_00_06 = i_multiplier[0] & i_multiplicand[6];
wire w_pp_00_07 = i_multiplier[0] & i_multiplicand[7];
wire w_pp_00_08 = i_multiplier[0] & i_multiplicand[8];
wire w_pp_00_09 = i_multiplier[0] & i_multiplicand[9];
wire w_pp_00_10 = i_multiplier[0] & i_multiplicand[10];
wire w_pp_00_11 = i_multiplier[0] & i_multiplicand[11];
wire w_pp_00_12 = i_multiplier[0] & i_multiplicand[12];
wire w_pp_00_13 = i_multiplier[0] & i_multiplicand[13];
wire w_pp_00_14 = i_multiplier[0] & i_multiplicand[14];
wire w_pp_00_15 = i_multiplier[0] & i_multiplicand[15];
wire w_pp_00_16 = i_multiplier[0] & i_multiplicand[16];
wire w_pp_00_17 = i_multiplier[0] & i_multiplicand[17];
wire w_pp_00_18 = i_multiplier[0] & i_multiplicand[18];
wire w_pp_00_19 = i_multiplier[0] & i_multiplicand[19];
wire w_pp_00_20 = i_multiplier[0] & i_multiplicand[20];
wire w_pp_00_21 = i_multiplier[0] & i_multiplicand[21];
wire w_pp_00_22 = i_multiplier[0] & i_multiplicand[22];
wire w_pp_00_23 = i_multiplier[0] & i_multiplicand[23];
wire w_pp_01_00 = i_multiplier[1] & i_multiplicand[0];
wire w_pp_01_01 = i_multiplier[1] & i_multiplicand[1];
wire w_pp_01_02 = i_multiplier[1] & i_multiplicand[2];
wire w_pp_01_03 = i_multiplier[1] & i_multiplicand[3];
wire w_pp_01_04 = i_multiplier[1] & i_multiplicand[4];
wire w_pp_01_05 = i_multiplier[1] & i_multiplicand[5];
wire w_pp_01_06 = i_multiplier[1] & i_multiplicand[6];
wire w_pp_01_07 = i_multiplier[1] & i_multiplicand[7];
wire w_pp_01_08 = i_multiplier[1] & i_multiplicand[8];
wire w_pp_01_09 = i_multiplier[1] & i_multiplicand[9];
wire w_pp_01_10 = i_multiplier[1] & i_multiplicand[10];
wire w_pp_01_11 = i_multiplier[1] & i_multiplicand[11];
wire w_pp_01_12 = i_multiplier[1] & i_multiplicand[12];
wire w_pp_01_13 = i_multiplier[1] & i_multiplicand[13];
wire w_pp_01_14 = i_multiplier[1] & i_multiplicand[14];
wire w_pp_01_15 = i_multiplier[1] & i_multiplicand[15];
wire w_pp_01_16 = i_multiplier[1] & i_multiplicand[16];
wire w_pp_01_17 = i_multiplier[1] & i_multiplicand[17];
wire w_pp_01_18 = i_multiplier[1] & i_multiplicand[18];
wire w_pp_01_19 = i_multiplier[1] & i_multiplicand[19];
wire w_pp_01_20 = i_multiplier[1] & i_multiplicand[20];
wire w_pp_01_21 = i_multiplier[1] & i_multiplicand[21];
wire w_pp_01_22 = i_multiplier[1] & i_multiplicand[22];
wire w_pp_01_23 = i_multiplier[1] & i_multiplicand[23];
wire w_pp_02_00 = i_multiplier[2] & i_multiplicand[0];
wire w_pp_02_01 = i_multiplier[2] & i_multiplicand[1];
wire w_pp_02_02 = i_multiplier[2] & i_multiplicand[2];
wire w_pp_02_03 = i_multiplier[2] & i_multiplicand[3];
wire w_pp_02_04 = i_multiplier[2] & i_multiplicand[4];
wire w_pp_02_05 = i_multiplier[2] & i_multiplicand[5];
wire w_pp_02_06 = i_multiplier[2] & i_multiplicand[6];
wire w_pp_02_07 = i_multiplier[2] & i_multiplicand[7];
wire w_pp_02_08 = i_multiplier[2] & i_multiplicand[8];
wire w_pp_02_09 = i_multiplier[2] & i_multiplicand[9];
wire w_pp_02_10 = i_multiplier[2] & i_multiplicand[10];
wire w_pp_02_11 = i_multiplier[2] & i_multiplicand[11];
wire w_pp_02_12 = i_multiplier[2] & i_multiplicand[12];
wire w_pp_02_13 = i_multiplier[2] & i_multiplicand[13];
wire w_pp_02_14 = i_multiplier[2] & i_multiplicand[14];
wire w_pp_02_15 = i_multiplier[2] & i_multiplicand[15];
wire w_pp_02_16 = i_multiplier[2] & i_multiplicand[16];
wire w_pp_02_17 = i_multiplier[2] & i_multiplicand[17];
wire w_pp_02_18 = i_multiplier[2] & i_multiplicand[18];
wire w_pp_02_19 = i_multiplier[2] & i_multiplicand[19];
wire w_pp_02_20 = i_multiplier[2] & i_multiplicand[20];
wire w_pp_02_21 = i_multiplier[2] & i_multiplicand[21];
wire w_pp_02_22 = i_multiplier[2] & i_multiplicand[22];
wire w_pp_02_23 = i_multiplier[2] & i_multiplicand[23];
wire w_pp_03_00 = i_multiplier[3] & i_multiplicand[0];
wire w_pp_03_01 = i_multiplier[3] & i_multiplicand[1];
wire w_pp_03_02 = i_multiplier[3] & i_multiplicand[2];
wire w_pp_03_03 = i_multiplier[3] & i_multiplicand[3];
wire w_pp_03_04 = i_multiplier[3] & i_multiplicand[4];
wire w_pp_03_05 = i_multiplier[3] & i_multiplicand[5];
wire w_pp_03_06 = i_multiplier[3] & i_multiplicand[6];
wire w_pp_03_07 = i_multiplier[3] & i_multiplicand[7];
wire w_pp_03_08 = i_multiplier[3] & i_multiplicand[8];
wire w_pp_03_09 = i_multiplier[3] & i_multiplicand[9];
wire w_pp_03_10 = i_multiplier[3] & i_multiplicand[10];
wire w_pp_03_11 = i_multiplier[3] & i_multiplicand[11];
wire w_pp_03_12 = i_multiplier[3] & i_multiplicand[12];
wire w_pp_03_13 = i_multiplier[3] & i_multiplicand[13];
wire w_pp_03_14 = i_multiplier[3] & i_multiplicand[14];
wire w_pp_03_15 = i_multiplier[3] & i_multiplicand[15];
wire w_pp_03_16 = i_multiplier[3] & i_multiplicand[16];
wire w_pp_03_17 = i_multiplier[3] & i_multiplicand[17];
wire w_pp_03_18 = i_multiplier[3] & i_multiplicand[18];
wire w_pp_03_19 = i_multiplier[3] & i_multiplicand[19];
wire w_pp_03_20 = i_multiplier[3] & i_multiplicand[20];
wire w_pp_03_21 = i_multiplier[3] & i_multiplicand[21];
wire w_pp_03_22 = i_multiplier[3] & i_multiplicand[22];
wire w_pp_03_23 = i_multiplier[3] & i_multiplicand[23];
wire w_pp_04_00 = i_multiplier[4] & i_multiplicand[0];
wire w_pp_04_01 = i_multiplier[4] & i_multiplicand[1];
wire w_pp_04_02 = i_multiplier[4] & i_multiplicand[2];
wire w_pp_04_03 = i_multiplier[4] & i_multiplicand[3];
wire w_pp_04_04 = i_multiplier[4] & i_multiplicand[4];
wire w_pp_04_05 = i_multiplier[4] & i_multiplicand[5];
wire w_pp_04_06 = i_multiplier[4] & i_multiplicand[6];
wire w_pp_04_07 = i_multiplier[4] & i_multiplicand[7];
wire w_pp_04_08 = i_multiplier[4] & i_multiplicand[8];
wire w_pp_04_09 = i_multiplier[4] & i_multiplicand[9];
wire w_pp_04_10 = i_multiplier[4] & i_multiplicand[10];
wire w_pp_04_11 = i_multiplier[4] & i_multiplicand[11];
wire w_pp_04_12 = i_multiplier[4] & i_multiplicand[12];
wire w_pp_04_13 = i_multiplier[4] & i_multiplicand[13];
wire w_pp_04_14 = i_multiplier[4] & i_multiplicand[14];
wire w_pp_04_15 = i_multiplier[4] & i_multiplicand[15];
wire w_pp_04_16 = i_multiplier[4] & i_multiplicand[16];
wire w_pp_04_17 = i_multiplier[4] & i_multiplicand[17];
wire w_pp_04_18 = i_multiplier[4] & i_multiplicand[18];
wire w_pp_04_19 = i_multiplier[4] & i_multiplicand[19];
wire w_pp_04_20 = i_multiplier[4] & i_multiplicand[20];
wire w_pp_04_21 = i_multiplier[4] & i_multiplicand[21];
wire w_pp_04_22 = i_multiplier[4] & i_multiplicand[22];
wire w_pp_04_23 = i_multiplier[4] & i_multiplicand[23];
wire w_pp_05_00 = i_multiplier[5] & i_multiplicand[0];
wire w_pp_05_01 = i_multiplier[5] & i_multiplicand[1];
wire w_pp_05_02 = i_multiplier[5] & i_multiplicand[2];
wire w_pp_05_03 = i_multiplier[5] & i_multiplicand[3];
wire w_pp_05_04 = i_multiplier[5] & i_multiplicand[4];
wire w_pp_05_05 = i_multiplier[5] & i_multiplicand[5];
wire w_pp_05_06 = i_multiplier[5] & i_multiplicand[6];
wire w_pp_05_07 = i_multiplier[5] & i_multiplicand[7];
wire w_pp_05_08 = i_multiplier[5] & i_multiplicand[8];
wire w_pp_05_09 = i_multiplier[5] & i_multiplicand[9];
wire w_pp_05_10 = i_multiplier[5] & i_multiplicand[10];
wire w_pp_05_11 = i_multiplier[5] & i_multiplicand[11];
wire w_pp_05_12 = i_multiplier[5] & i_multiplicand[12];
wire w_pp_05_13 = i_multiplier[5] & i_multiplicand[13];
wire w_pp_05_14 = i_multiplier[5] & i_multiplicand[14];
wire w_pp_05_15 = i_multiplier[5] & i_multiplicand[15];
wire w_pp_05_16 = i_multiplier[5] & i_multiplicand[16];
wire w_pp_05_17 = i_multiplier[5] & i_multiplicand[17];
wire w_pp_05_18 = i_multiplier[5] & i_multiplicand[18];
wire w_pp_05_19 = i_multiplier[5] & i_multiplicand[19];
wire w_pp_05_20 = i_multiplier[5] & i_multiplicand[20];
wire w_pp_05_21 = i_multiplier[5] & i_multiplicand[21];
wire w_pp_05_22 = i_multiplier[5] & i_multiplicand[22];
wire w_pp_05_23 = i_multiplier[5] & i_multiplicand[23];
wire w_pp_06_00 = i_multiplier[6] & i_multiplicand[0];
wire w_pp_06_01 = i_multiplier[6] & i_multiplicand[1];
wire w_pp_06_02 = i_multiplier[6] & i_multiplicand[2];
wire w_pp_06_03 = i_multiplier[6] & i_multiplicand[3];
wire w_pp_06_04 = i_multiplier[6] & i_multiplicand[4];
wire w_pp_06_05 = i_multiplier[6] & i_multiplicand[5];
wire w_pp_06_06 = i_multiplier[6] & i_multiplicand[6];
wire w_pp_06_07 = i_multiplier[6] & i_multiplicand[7];
wire w_pp_06_08 = i_multiplier[6] & i_multiplicand[8];
wire w_pp_06_09 = i_multiplier[6] & i_multiplicand[9];
wire w_pp_06_10 = i_multiplier[6] & i_multiplicand[10];
wire w_pp_06_11 = i_multiplier[6] & i_multiplicand[11];
wire w_pp_06_12 = i_multiplier[6] & i_multiplicand[12];
wire w_pp_06_13 = i_multiplier[6] & i_multiplicand[13];
wire w_pp_06_14 = i_multiplier[6] & i_multiplicand[14];
wire w_pp_06_15 = i_multiplier[6] & i_multiplicand[15];
wire w_pp_06_16 = i_multiplier[6] & i_multiplicand[16];
wire w_pp_06_17 = i_multiplier[6] & i_multiplicand[17];
wire w_pp_06_18 = i_multiplier[6] & i_multiplicand[18];
wire w_pp_06_19 = i_multiplier[6] & i_multiplicand[19];
wire w_pp_06_20 = i_multiplier[6] & i_multiplicand[20];
wire w_pp_06_21 = i_multiplier[6] & i_multiplicand[21];
wire w_pp_06_22 = i_multiplier[6] & i_multiplicand[22];
wire w_pp_06_23 = i_multiplier[6] & i_multiplicand[23];
wire w_pp_07_00 = i_multiplier[7] & i_multiplicand[0];
wire w_pp_07_01 = i_multiplier[7] & i_multiplicand[1];
wire w_pp_07_02 = i_multiplier[7] & i_multiplicand[2];
wire w_pp_07_03 = i_multiplier[7] & i_multiplicand[3];
wire w_pp_07_04 = i_multiplier[7] & i_multiplicand[4];
wire w_pp_07_05 = i_multiplier[7] & i_multiplicand[5];
wire w_pp_07_06 = i_multiplier[7] & i_multiplicand[6];
wire w_pp_07_07 = i_multiplier[7] & i_multiplicand[7];
wire w_pp_07_08 = i_multiplier[7] & i_multiplicand[8];
wire w_pp_07_09 = i_multiplier[7] & i_multiplicand[9];
wire w_pp_07_10 = i_multiplier[7] & i_multiplicand[10];
wire w_pp_07_11 = i_multiplier[7] & i_multiplicand[11];
wire w_pp_07_12 = i_multiplier[7] & i_multiplicand[12];
wire w_pp_07_13 = i_multiplier[7] & i_multiplicand[13];
wire w_pp_07_14 = i_multiplier[7] & i_multiplicand[14];
wire w_pp_07_15 = i_multiplier[7] & i_multiplicand[15];
wire w_pp_07_16 = i_multiplier[7] & i_multiplicand[16];
wire w_pp_07_17 = i_multiplier[7] & i_multiplicand[17];
wire w_pp_07_18 = i_multiplier[7] & i_multiplicand[18];
wire w_pp_07_19 = i_multiplier[7] & i_multiplicand[19];
wire w_pp_07_20 = i_multiplier[7] & i_multiplicand[20];
wire w_pp_07_21 = i_multiplier[7] & i_multiplicand[21];
wire w_pp_07_22 = i_multiplier[7] & i_multiplicand[22];
wire w_pp_07_23 = i_multiplier[7] & i_multiplicand[23];
wire w_pp_08_00 = i_multiplier[8] & i_multiplicand[0];
wire w_pp_08_01 = i_multiplier[8] & i_multiplicand[1];
wire w_pp_08_02 = i_multiplier[8] & i_multiplicand[2];
wire w_pp_08_03 = i_multiplier[8] & i_multiplicand[3];
wire w_pp_08_04 = i_multiplier[8] & i_multiplicand[4];
wire w_pp_08_05 = i_multiplier[8] & i_multiplicand[5];
wire w_pp_08_06 = i_multiplier[8] & i_multiplicand[6];
wire w_pp_08_07 = i_multiplier[8] & i_multiplicand[7];
wire w_pp_08_08 = i_multiplier[8] & i_multiplicand[8];
wire w_pp_08_09 = i_multiplier[8] & i_multiplicand[9];
wire w_pp_08_10 = i_multiplier[8] & i_multiplicand[10];
wire w_pp_08_11 = i_multiplier[8] & i_multiplicand[11];
wire w_pp_08_12 = i_multiplier[8] & i_multiplicand[12];
wire w_pp_08_13 = i_multiplier[8] & i_multiplicand[13];
wire w_pp_08_14 = i_multiplier[8] & i_multiplicand[14];
wire w_pp_08_15 = i_multiplier[8] & i_multiplicand[15];
wire w_pp_08_16 = i_multiplier[8] & i_multiplicand[16];
wire w_pp_08_17 = i_multiplier[8] & i_multiplicand[17];
wire w_pp_08_18 = i_multiplier[8] & i_multiplicand[18];
wire w_pp_08_19 = i_multiplier[8] & i_multiplicand[19];
wire w_pp_08_20 = i_multiplier[8] & i_multiplicand[20];
wire w_pp_08_21 = i_multiplier[8] & i_multiplicand[21];
wire w_pp_08_22 = i_multiplier[8] & i_multiplicand[22];
wire w_pp_08_23 = i_multiplier[8] & i_multiplicand[23];
wire w_pp_09_00 = i_multiplier[9] & i_multiplicand[0];
wire w_pp_09_01 = i_multiplier[9] & i_multiplicand[1];
wire w_pp_09_02 = i_multiplier[9] & i_multiplicand[2];
wire w_pp_09_03 = i_multiplier[9] & i_multiplicand[3];
wire w_pp_09_04 = i_multiplier[9] & i_multiplicand[4];
wire w_pp_09_05 = i_multiplier[9] & i_multiplicand[5];
wire w_pp_09_06 = i_multiplier[9] & i_multiplicand[6];
wire w_pp_09_07 = i_multiplier[9] & i_multiplicand[7];
wire w_pp_09_08 = i_multiplier[9] & i_multiplicand[8];
wire w_pp_09_09 = i_multiplier[9] & i_multiplicand[9];
wire w_pp_09_10 = i_multiplier[9] & i_multiplicand[10];
wire w_pp_09_11 = i_multiplier[9] & i_multiplicand[11];
wire w_pp_09_12 = i_multiplier[9] & i_multiplicand[12];
wire w_pp_09_13 = i_multiplier[9] & i_multiplicand[13];
wire w_pp_09_14 = i_multiplier[9] & i_multiplicand[14];
wire w_pp_09_15 = i_multiplier[9] & i_multiplicand[15];
wire w_pp_09_16 = i_multiplier[9] & i_multiplicand[16];
wire w_pp_09_17 = i_multiplier[9] & i_multiplicand[17];
wire w_pp_09_18 = i_multiplier[9] & i_multiplicand[18];
wire w_pp_09_19 = i_multiplier[9] & i_multiplicand[19];
wire w_pp_09_20 = i_multiplier[9] & i_multiplicand[20];
wire w_pp_09_21 = i_multiplier[9] & i_multiplicand[21];
wire w_pp_09_22 = i_multiplier[9] & i_multiplicand[22];
wire w_pp_09_23 = i_multiplier[9] & i_multiplicand[23];
wire w_pp_10_00 = i_multiplier[10] & i_multiplicand[0];
wire w_pp_10_01 = i_multiplier[10] & i_multiplicand[1];
wire w_pp_10_02 = i_multiplier[10] & i_multiplicand[2];
wire w_pp_10_03 = i_multiplier[10] & i_multiplicand[3];
wire w_pp_10_04 = i_multiplier[10] & i_multiplicand[4];
wire w_pp_10_05 = i_multiplier[10] & i_multiplicand[5];
wire w_pp_10_06 = i_multiplier[10] & i_multiplicand[6];
wire w_pp_10_07 = i_multiplier[10] & i_multiplicand[7];
wire w_pp_10_08 = i_multiplier[10] & i_multiplicand[8];
wire w_pp_10_09 = i_multiplier[10] & i_multiplicand[9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_10_16 = i_multiplier[10] & i_multiplicand[16];
wire w_pp_10_17 = i_multiplier[10] & i_multiplicand[17];
wire w_pp_10_18 = i_multiplier[10] & i_multiplicand[18];
wire w_pp_10_19 = i_multiplier[10] & i_multiplicand[19];
wire w_pp_10_20 = i_multiplier[10] & i_multiplicand[20];
wire w_pp_10_21 = i_multiplier[10] & i_multiplicand[21];
wire w_pp_10_22 = i_multiplier[10] & i_multiplicand[22];
wire w_pp_10_23 = i_multiplier[10] & i_multiplicand[23];
wire w_pp_11_00 = i_multiplier[11] & i_multiplicand[0];
wire w_pp_11_01 = i_multiplier[11] & i_multiplicand[1];
wire w_pp_11_02 = i_multiplier[11] & i_multiplicand[2];
wire w_pp_11_03 = i_multiplier[11] & i_multiplicand[3];
wire w_pp_11_04 = i_multiplier[11] & i_multiplicand[4];
wire w_pp_11_05 = i_multiplier[11] & i_multiplicand[5];
wire w_pp_11_06 = i_multiplier[11] & i_multiplicand[6];
wire w_pp_11_07 = i_multiplier[11] & i_multiplicand[7];
wire w_pp_11_08 = i_multiplier[11] & i_multiplicand[8];
wire w_pp_11_09 = i_multiplier[11] & i_multiplicand[9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_11_16 = i_multiplier[11] & i_multiplicand[16];
wire w_pp_11_17 = i_multiplier[11] & i_multiplicand[17];
wire w_pp_11_18 = i_multiplier[11] & i_multiplicand[18];
wire w_pp_11_19 = i_multiplier[11] & i_multiplicand[19];
wire w_pp_11_20 = i_multiplier[11] & i_multiplicand[20];
wire w_pp_11_21 = i_multiplier[11] & i_multiplicand[21];
wire w_pp_11_22 = i_multiplier[11] & i_multiplicand[22];
wire w_pp_11_23 = i_multiplier[11] & i_multiplicand[23];
wire w_pp_12_00 = i_multiplier[12] & i_multiplicand[0];
wire w_pp_12_01 = i_multiplier[12] & i_multiplicand[1];
wire w_pp_12_02 = i_multiplier[12] & i_multiplicand[2];
wire w_pp_12_03 = i_multiplier[12] & i_multiplicand[3];
wire w_pp_12_04 = i_multiplier[12] & i_multiplicand[4];
wire w_pp_12_05 = i_multiplier[12] & i_multiplicand[5];
wire w_pp_12_06 = i_multiplier[12] & i_multiplicand[6];
wire w_pp_12_07 = i_multiplier[12] & i_multiplicand[7];
wire w_pp_12_08 = i_multiplier[12] & i_multiplicand[8];
wire w_pp_12_09 = i_multiplier[12] & i_multiplicand[9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_12_16 = i_multiplier[12] & i_multiplicand[16];
wire w_pp_12_17 = i_multiplier[12] & i_multiplicand[17];
wire w_pp_12_18 = i_multiplier[12] & i_multiplicand[18];
wire w_pp_12_19 = i_multiplier[12] & i_multiplicand[19];
wire w_pp_12_20 = i_multiplier[12] & i_multiplicand[20];
wire w_pp_12_21 = i_multiplier[12] & i_multiplicand[21];
wire w_pp_12_22 = i_multiplier[12] & i_multiplicand[22];
wire w_pp_12_23 = i_multiplier[12] & i_multiplicand[23];
wire w_pp_13_00 = i_multiplier[13] & i_multiplicand[0];
wire w_pp_13_01 = i_multiplier[13] & i_multiplicand[1];
wire w_pp_13_02 = i_multiplier[13] & i_multiplicand[2];
wire w_pp_13_03 = i_multiplier[13] & i_multiplicand[3];
wire w_pp_13_04 = i_multiplier[13] & i_multiplicand[4];
wire w_pp_13_05 = i_multiplier[13] & i_multiplicand[5];
wire w_pp_13_06 = i_multiplier[13] & i_multiplicand[6];
wire w_pp_13_07 = i_multiplier[13] & i_multiplicand[7];
wire w_pp_13_08 = i_multiplier[13] & i_multiplicand[8];
wire w_pp_13_09 = i_multiplier[13] & i_multiplicand[9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_13_16 = i_multiplier[13] & i_multiplicand[16];
wire w_pp_13_17 = i_multiplier[13] & i_multiplicand[17];
wire w_pp_13_18 = i_multiplier[13] & i_multiplicand[18];
wire w_pp_13_19 = i_multiplier[13] & i_multiplicand[19];
wire w_pp_13_20 = i_multiplier[13] & i_multiplicand[20];
wire w_pp_13_21 = i_multiplier[13] & i_multiplicand[21];
wire w_pp_13_22 = i_multiplier[13] & i_multiplicand[22];
wire w_pp_13_23 = i_multiplier[13] & i_multiplicand[23];
wire w_pp_14_00 = i_multiplier[14] & i_multiplicand[0];
wire w_pp_14_01 = i_multiplier[14] & i_multiplicand[1];
wire w_pp_14_02 = i_multiplier[14] & i_multiplicand[2];
wire w_pp_14_03 = i_multiplier[14] & i_multiplicand[3];
wire w_pp_14_04 = i_multiplier[14] & i_multiplicand[4];
wire w_pp_14_05 = i_multiplier[14] & i_multiplicand[5];
wire w_pp_14_06 = i_multiplier[14] & i_multiplicand[6];
wire w_pp_14_07 = i_multiplier[14] & i_multiplicand[7];
wire w_pp_14_08 = i_multiplier[14] & i_multiplicand[8];
wire w_pp_14_09 = i_multiplier[14] & i_multiplicand[9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_14_16 = i_multiplier[14] & i_multiplicand[16];
wire w_pp_14_17 = i_multiplier[14] & i_multiplicand[17];
wire w_pp_14_18 = i_multiplier[14] & i_multiplicand[18];
wire w_pp_14_19 = i_multiplier[14] & i_multiplicand[19];
wire w_pp_14_20 = i_multiplier[14] & i_multiplicand[20];
wire w_pp_14_21 = i_multiplier[14] & i_multiplicand[21];
wire w_pp_14_22 = i_multiplier[14] & i_multiplicand[22];
wire w_pp_14_23 = i_multiplier[14] & i_multiplicand[23];
wire w_pp_15_00 = i_multiplier[15] & i_multiplicand[0];
wire w_pp_15_01 = i_multiplier[15] & i_multiplicand[1];
wire w_pp_15_02 = i_multiplier[15] & i_multiplicand[2];
wire w_pp_15_03 = i_multiplier[15] & i_multiplicand[3];
wire w_pp_15_04 = i_multiplier[15] & i_multiplicand[4];
wire w_pp_15_05 = i_multiplier[15] & i_multiplicand[5];
wire w_pp_15_06 = i_multiplier[15] & i_multiplicand[6];
wire w_pp_15_07 = i_multiplier[15] & i_multiplicand[7];
wire w_pp_15_08 = i_multiplier[15] & i_multiplicand[8];
wire w_pp_15_09 = i_multiplier[15] & i_multiplicand[9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];
wire w_pp_15_16 = i_multiplier[15] & i_multiplicand[16];
wire w_pp_15_17 = i_multiplier[15] & i_multiplicand[17];
wire w_pp_15_18 = i_multiplier[15] & i_multiplicand[18];
wire w_pp_15_19 = i_multiplier[15] & i_multiplicand[19];
wire w_pp_15_20 = i_multiplier[15] & i_multiplicand[20];
wire w_pp_15_21 = i_multiplier[15] & i_multiplicand[21];
wire w_pp_15_22 = i_multiplier[15] & i_multiplicand[22];
wire w_pp_15_23 = i_multiplier[15] & i_multiplicand[23];
wire w_pp_16_00 = i_multiplier[16] & i_multiplicand[0];
wire w_pp_16_01 = i_multiplier[16] & i_multiplicand[1];
wire w_pp_16_02 = i_multiplier[16] & i_multiplicand[2];
wire w_pp_16_03 = i_multiplier[16] & i_multiplicand[3];
wire w_pp_16_04 = i_multiplier[16] & i_multiplicand[4];
wire w_pp_16_05 = i_multiplier[16] & i_multiplicand[5];
wire w_pp_16_06 = i_multiplier[16] & i_multiplicand[6];
wire w_pp_16_07 = i_multiplier[16] & i_multiplicand[7];
wire w_pp_16_08 = i_multiplier[16] & i_multiplicand[8];
wire w_pp_16_09 = i_multiplier[16] & i_multiplicand[9];
wire w_pp_16_10 = i_multiplier[16] & i_multiplicand[10];
wire w_pp_16_11 = i_multiplier[16] & i_multiplicand[11];
wire w_pp_16_12 = i_multiplier[16] & i_multiplicand[12];
wire w_pp_16_13 = i_multiplier[16] & i_multiplicand[13];
wire w_pp_16_14 = i_multiplier[16] & i_multiplicand[14];
wire w_pp_16_15 = i_multiplier[16] & i_multiplicand[15];
wire w_pp_16_16 = i_multiplier[16] & i_multiplicand[16];
wire w_pp_16_17 = i_multiplier[16] & i_multiplicand[17];
wire w_pp_16_18 = i_multiplier[16] & i_multiplicand[18];
wire w_pp_16_19 = i_multiplier[16] & i_multiplicand[19];
wire w_pp_16_20 = i_multiplier[16] & i_multiplicand[20];
wire w_pp_16_21 = i_multiplier[16] & i_multiplicand[21];
wire w_pp_16_22 = i_multiplier[16] & i_multiplicand[22];
wire w_pp_16_23 = i_multiplier[16] & i_multiplicand[23];
wire w_pp_17_00 = i_multiplier[17] & i_multiplicand[0];
wire w_pp_17_01 = i_multiplier[17] & i_multiplicand[1];
wire w_pp_17_02 = i_multiplier[17] & i_multiplicand[2];
wire w_pp_17_03 = i_multiplier[17] & i_multiplicand[3];
wire w_pp_17_04 = i_multiplier[17] & i_multiplicand[4];
wire w_pp_17_05 = i_multiplier[17] & i_multiplicand[5];
wire w_pp_17_06 = i_multiplier[17] & i_multiplicand[6];
wire w_pp_17_07 = i_multiplier[17] & i_multiplicand[7];
wire w_pp_17_08 = i_multiplier[17] & i_multiplicand[8];
wire w_pp_17_09 = i_multiplier[17] & i_multiplicand[9];
wire w_pp_17_10 = i_multiplier[17] & i_multiplicand[10];
wire w_pp_17_11 = i_multiplier[17] & i_multiplicand[11];
wire w_pp_17_12 = i_multiplier[17] & i_multiplicand[12];
wire w_pp_17_13 = i_multiplier[17] & i_multiplicand[13];
wire w_pp_17_14 = i_multiplier[17] & i_multiplicand[14];
wire w_pp_17_15 = i_multiplier[17] & i_multiplicand[15];
wire w_pp_17_16 = i_multiplier[17] & i_multiplicand[16];
wire w_pp_17_17 = i_multiplier[17] & i_multiplicand[17];
wire w_pp_17_18 = i_multiplier[17] & i_multiplicand[18];
wire w_pp_17_19 = i_multiplier[17] & i_multiplicand[19];
wire w_pp_17_20 = i_multiplier[17] & i_multiplicand[20];
wire w_pp_17_21 = i_multiplier[17] & i_multiplicand[21];
wire w_pp_17_22 = i_multiplier[17] & i_multiplicand[22];
wire w_pp_17_23 = i_multiplier[17] & i_multiplicand[23];
wire w_pp_18_00 = i_multiplier[18] & i_multiplicand[0];
wire w_pp_18_01 = i_multiplier[18] & i_multiplicand[1];
wire w_pp_18_02 = i_multiplier[18] & i_multiplicand[2];
wire w_pp_18_03 = i_multiplier[18] & i_multiplicand[3];
wire w_pp_18_04 = i_multiplier[18] & i_multiplicand[4];
wire w_pp_18_05 = i_multiplier[18] & i_multiplicand[5];
wire w_pp_18_06 = i_multiplier[18] & i_multiplicand[6];
wire w_pp_18_07 = i_multiplier[18] & i_multiplicand[7];
wire w_pp_18_08 = i_multiplier[18] & i_multiplicand[8];
wire w_pp_18_09 = i_multiplier[18] & i_multiplicand[9];
wire w_pp_18_10 = i_multiplier[18] & i_multiplicand[10];
wire w_pp_18_11 = i_multiplier[18] & i_multiplicand[11];
wire w_pp_18_12 = i_multiplier[18] & i_multiplicand[12];
wire w_pp_18_13 = i_multiplier[18] & i_multiplicand[13];
wire w_pp_18_14 = i_multiplier[18] & i_multiplicand[14];
wire w_pp_18_15 = i_multiplier[18] & i_multiplicand[15];
wire w_pp_18_16 = i_multiplier[18] & i_multiplicand[16];
wire w_pp_18_17 = i_multiplier[18] & i_multiplicand[17];
wire w_pp_18_18 = i_multiplier[18] & i_multiplicand[18];
wire w_pp_18_19 = i_multiplier[18] & i_multiplicand[19];
wire w_pp_18_20 = i_multiplier[18] & i_multiplicand[20];
wire w_pp_18_21 = i_multiplier[18] & i_multiplicand[21];
wire w_pp_18_22 = i_multiplier[18] & i_multiplicand[22];
wire w_pp_18_23 = i_multiplier[18] & i_multiplicand[23];
wire w_pp_19_00 = i_multiplier[19] & i_multiplicand[0];
wire w_pp_19_01 = i_multiplier[19] & i_multiplicand[1];
wire w_pp_19_02 = i_multiplier[19] & i_multiplicand[2];
wire w_pp_19_03 = i_multiplier[19] & i_multiplicand[3];
wire w_pp_19_04 = i_multiplier[19] & i_multiplicand[4];
wire w_pp_19_05 = i_multiplier[19] & i_multiplicand[5];
wire w_pp_19_06 = i_multiplier[19] & i_multiplicand[6];
wire w_pp_19_07 = i_multiplier[19] & i_multiplicand[7];
wire w_pp_19_08 = i_multiplier[19] & i_multiplicand[8];
wire w_pp_19_09 = i_multiplier[19] & i_multiplicand[9];
wire w_pp_19_10 = i_multiplier[19] & i_multiplicand[10];
wire w_pp_19_11 = i_multiplier[19] & i_multiplicand[11];
wire w_pp_19_12 = i_multiplier[19] & i_multiplicand[12];
wire w_pp_19_13 = i_multiplier[19] & i_multiplicand[13];
wire w_pp_19_14 = i_multiplier[19] & i_multiplicand[14];
wire w_pp_19_15 = i_multiplier[19] & i_multiplicand[15];
wire w_pp_19_16 = i_multiplier[19] & i_multiplicand[16];
wire w_pp_19_17 = i_multiplier[19] & i_multiplicand[17];
wire w_pp_19_18 = i_multiplier[19] & i_multiplicand[18];
wire w_pp_19_19 = i_multiplier[19] & i_multiplicand[19];
wire w_pp_19_20 = i_multiplier[19] & i_multiplicand[20];
wire w_pp_19_21 = i_multiplier[19] & i_multiplicand[21];
wire w_pp_19_22 = i_multiplier[19] & i_multiplicand[22];
wire w_pp_19_23 = i_multiplier[19] & i_multiplicand[23];
wire w_pp_20_00 = i_multiplier[20] & i_multiplicand[0];
wire w_pp_20_01 = i_multiplier[20] & i_multiplicand[1];
wire w_pp_20_02 = i_multiplier[20] & i_multiplicand[2];
wire w_pp_20_03 = i_multiplier[20] & i_multiplicand[3];
wire w_pp_20_04 = i_multiplier[20] & i_multiplicand[4];
wire w_pp_20_05 = i_multiplier[20] & i_multiplicand[5];
wire w_pp_20_06 = i_multiplier[20] & i_multiplicand[6];
wire w_pp_20_07 = i_multiplier[20] & i_multiplicand[7];
wire w_pp_20_08 = i_multiplier[20] & i_multiplicand[8];
wire w_pp_20_09 = i_multiplier[20] & i_multiplicand[9];
wire w_pp_20_10 = i_multiplier[20] & i_multiplicand[10];
wire w_pp_20_11 = i_multiplier[20] & i_multiplicand[11];
wire w_pp_20_12 = i_multiplier[20] & i_multiplicand[12];
wire w_pp_20_13 = i_multiplier[20] & i_multiplicand[13];
wire w_pp_20_14 = i_multiplier[20] & i_multiplicand[14];
wire w_pp_20_15 = i_multiplier[20] & i_multiplicand[15];
wire w_pp_20_16 = i_multiplier[20] & i_multiplicand[16];
wire w_pp_20_17 = i_multiplier[20] & i_multiplicand[17];
wire w_pp_20_18 = i_multiplier[20] & i_multiplicand[18];
wire w_pp_20_19 = i_multiplier[20] & i_multiplicand[19];
wire w_pp_20_20 = i_multiplier[20] & i_multiplicand[20];
wire w_pp_20_21 = i_multiplier[20] & i_multiplicand[21];
wire w_pp_20_22 = i_multiplier[20] & i_multiplicand[22];
wire w_pp_20_23 = i_multiplier[20] & i_multiplicand[23];
wire w_pp_21_00 = i_multiplier[21] & i_multiplicand[0];
wire w_pp_21_01 = i_multiplier[21] & i_multiplicand[1];
wire w_pp_21_02 = i_multiplier[21] & i_multiplicand[2];
wire w_pp_21_03 = i_multiplier[21] & i_multiplicand[3];
wire w_pp_21_04 = i_multiplier[21] & i_multiplicand[4];
wire w_pp_21_05 = i_multiplier[21] & i_multiplicand[5];
wire w_pp_21_06 = i_multiplier[21] & i_multiplicand[6];
wire w_pp_21_07 = i_multiplier[21] & i_multiplicand[7];
wire w_pp_21_08 = i_multiplier[21] & i_multiplicand[8];
wire w_pp_21_09 = i_multiplier[21] & i_multiplicand[9];
wire w_pp_21_10 = i_multiplier[21] & i_multiplicand[10];
wire w_pp_21_11 = i_multiplier[21] & i_multiplicand[11];
wire w_pp_21_12 = i_multiplier[21] & i_multiplicand[12];
wire w_pp_21_13 = i_multiplier[21] & i_multiplicand[13];
wire w_pp_21_14 = i_multiplier[21] & i_multiplicand[14];
wire w_pp_21_15 = i_multiplier[21] & i_multiplicand[15];
wire w_pp_21_16 = i_multiplier[21] & i_multiplicand[16];
wire w_pp_21_17 = i_multiplier[21] & i_multiplicand[17];
wire w_pp_21_18 = i_multiplier[21] & i_multiplicand[18];
wire w_pp_21_19 = i_multiplier[21] & i_multiplicand[19];
wire w_pp_21_20 = i_multiplier[21] & i_multiplicand[20];
wire w_pp_21_21 = i_multiplier[21] & i_multiplicand[21];
wire w_pp_21_22 = i_multiplier[21] & i_multiplicand[22];
wire w_pp_21_23 = i_multiplier[21] & i_multiplicand[23];
wire w_pp_22_00 = i_multiplier[22] & i_multiplicand[0];
wire w_pp_22_01 = i_multiplier[22] & i_multiplicand[1];
wire w_pp_22_02 = i_multiplier[22] & i_multiplicand[2];
wire w_pp_22_03 = i_multiplier[22] & i_multiplicand[3];
wire w_pp_22_04 = i_multiplier[22] & i_multiplicand[4];
wire w_pp_22_05 = i_multiplier[22] & i_multiplicand[5];
wire w_pp_22_06 = i_multiplier[22] & i_multiplicand[6];
wire w_pp_22_07 = i_multiplier[22] & i_multiplicand[7];
wire w_pp_22_08 = i_multiplier[22] & i_multiplicand[8];
wire w_pp_22_09 = i_multiplier[22] & i_multiplicand[9];
wire w_pp_22_10 = i_multiplier[22] & i_multiplicand[10];
wire w_pp_22_11 = i_multiplier[22] & i_multiplicand[11];
wire w_pp_22_12 = i_multiplier[22] & i_multiplicand[12];
wire w_pp_22_13 = i_multiplier[22] & i_multiplicand[13];
wire w_pp_22_14 = i_multiplier[22] & i_multiplicand[14];
wire w_pp_22_15 = i_multiplier[22] & i_multiplicand[15];
wire w_pp_22_16 = i_multiplier[22] & i_multiplicand[16];
wire w_pp_22_17 = i_multiplier[22] & i_multiplicand[17];
wire w_pp_22_18 = i_multiplier[22] & i_multiplicand[18];
wire w_pp_22_19 = i_multiplier[22] & i_multiplicand[19];
wire w_pp_22_20 = i_multiplier[22] & i_multiplicand[20];
wire w_pp_22_21 = i_multiplier[22] & i_multiplicand[21];
wire w_pp_22_22 = i_multiplier[22] & i_multiplicand[22];
wire w_pp_22_23 = i_multiplier[22] & i_multiplicand[23];
wire w_pp_23_00 = i_multiplier[23] & i_multiplicand[0];
wire w_pp_23_01 = i_multiplier[23] & i_multiplicand[1];
wire w_pp_23_02 = i_multiplier[23] & i_multiplicand[2];
wire w_pp_23_03 = i_multiplier[23] & i_multiplicand[3];
wire w_pp_23_04 = i_multiplier[23] & i_multiplicand[4];
wire w_pp_23_05 = i_multiplier[23] & i_multiplicand[5];
wire w_pp_23_06 = i_multiplier[23] & i_multiplicand[6];
wire w_pp_23_07 = i_multiplier[23] & i_multiplicand[7];
wire w_pp_23_08 = i_multiplier[23] & i_multiplicand[8];
wire w_pp_23_09 = i_multiplier[23] & i_multiplicand[9];
wire w_pp_23_10 = i_multiplier[23] & i_multiplicand[10];
wire w_pp_23_11 = i_multiplier[23] & i_multiplicand[11];
wire w_pp_23_12 = i_multiplier[23] & i_multiplicand[12];
wire w_pp_23_13 = i_multiplier[23] & i_multiplicand[13];
wire w_pp_23_14 = i_multiplier[23] & i_multiplicand[14];
wire w_pp_23_15 = i_multiplier[23] & i_multiplicand[15];
wire w_pp_23_16 = i_multiplier[23] & i_multiplicand[16];
wire w_pp_23_17 = i_multiplier[23] & i_multiplicand[17];
wire w_pp_23_18 = i_multiplier[23] & i_multiplicand[18];
wire w_pp_23_19 = i_multiplier[23] & i_multiplicand[19];
wire w_pp_23_20 = i_multiplier[23] & i_multiplicand[20];
wire w_pp_23_21 = i_multiplier[23] & i_multiplicand[21];
wire w_pp_23_22 = i_multiplier[23] & i_multiplicand[22];
wire w_pp_23_23 = i_multiplier[23] & i_multiplicand[23];

// Dadda Reduction Stage 1: height 24 -> 19

wire w_c4to2_sum_19_000, w_c4to2_carry_19_000, w_c4to2_cout_19_000;
math_compressor_4to2 u_c4to2_19_000 (
    .i_x1(w_pp_00_19), .i_x2(w_pp_01_18),
    .i_x3(w_pp_02_17), .i_x4(w_pp_03_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_000), .ow_carry(w_c4to2_carry_19_000), .ow_cout(w_c4to2_cout_19_000)
);
wire w_c4to2_sum_20_001, w_c4to2_carry_20_001, w_c4to2_cout_20_001;
math_compressor_4to2 u_c4to2_20_001 (
    .i_x1(w_pp_00_20), .i_x2(w_pp_01_19),
    .i_x3(w_pp_02_18), .i_x4(w_pp_03_17),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_001), .ow_carry(w_c4to2_carry_20_001), .ow_cout(w_c4to2_cout_20_001)
);
wire w_c4to2_sum_20_002, w_c4to2_carry_20_002, w_c4to2_cout_20_002;
math_compressor_4to2 u_c4to2_20_002 (
    .i_x1(w_pp_04_16), .i_x2(w_pp_05_15),
    .i_x3(w_pp_06_14), .i_x4(w_pp_07_13),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_002), .ow_carry(w_c4to2_carry_20_002), .ow_cout(w_c4to2_cout_20_002)
);
wire w_c4to2_sum_21_003, w_c4to2_carry_21_003, w_c4to2_cout_21_003;
math_compressor_4to2 u_c4to2_21_003 (
    .i_x1(w_pp_00_21), .i_x2(w_pp_01_20),
    .i_x3(w_pp_02_19), .i_x4(w_pp_03_18),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_003), .ow_carry(w_c4to2_carry_21_003), .ow_cout(w_c4to2_cout_21_003)
);
wire w_c4to2_sum_21_004, w_c4to2_carry_21_004, w_c4to2_cout_21_004;
math_compressor_4to2 u_c4to2_21_004 (
    .i_x1(w_pp_04_17), .i_x2(w_pp_05_16),
    .i_x3(w_pp_06_15), .i_x4(w_pp_07_14),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_004), .ow_carry(w_c4to2_carry_21_004), .ow_cout(w_c4to2_cout_21_004)
);
wire w_c4to2_sum_21_005, w_c4to2_carry_21_005, w_c4to2_cout_21_005;
math_compressor_4to2 u_c4to2_21_005 (
    .i_x1(w_pp_08_13), .i_x2(w_pp_09_12),
    .i_x3(w_pp_10_11), .i_x4(w_pp_11_10),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_005), .ow_carry(w_c4to2_carry_21_005), .ow_cout(w_c4to2_cout_21_005)
);
wire w_c4to2_sum_22_006, w_c4to2_carry_22_006, w_c4to2_cout_22_006;
math_compressor_4to2 u_c4to2_22_006 (
    .i_x1(w_pp_00_22), .i_x2(w_pp_01_21),
    .i_x3(w_pp_02_20), .i_x4(w_pp_03_19),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_006), .ow_carry(w_c4to2_carry_22_006), .ow_cout(w_c4to2_cout_22_006)
);
wire w_c4to2_sum_22_007, w_c4to2_carry_22_007, w_c4to2_cout_22_007;
math_compressor_4to2 u_c4to2_22_007 (
    .i_x1(w_pp_04_18), .i_x2(w_pp_05_17),
    .i_x3(w_pp_06_16), .i_x4(w_pp_07_15),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_007), .ow_carry(w_c4to2_carry_22_007), .ow_cout(w_c4to2_cout_22_007)
);
wire w_c4to2_sum_22_008, w_c4to2_carry_22_008, w_c4to2_cout_22_008;
math_compressor_4to2 u_c4to2_22_008 (
    .i_x1(w_pp_08_14), .i_x2(w_pp_09_13),
    .i_x3(w_pp_10_12), .i_x4(w_pp_11_11),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_008), .ow_carry(w_c4to2_carry_22_008), .ow_cout(w_c4to2_cout_22_008)
);
wire w_c4to2_sum_22_009, w_c4to2_carry_22_009, w_c4to2_cout_22_009;
math_compressor_4to2 u_c4to2_22_009 (
    .i_x1(w_pp_12_10), .i_x2(w_pp_13_09),
    .i_x3(w_pp_14_08), .i_x4(w_pp_15_07),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_009), .ow_carry(w_c4to2_carry_22_009), .ow_cout(w_c4to2_cout_22_009)
);
wire w_c4to2_sum_23_010, w_c4to2_carry_23_010, w_c4to2_cout_23_010;
math_compressor_4to2 u_c4to2_23_010 (
    .i_x1(w_pp_00_23), .i_x2(w_pp_01_22),
    .i_x3(w_pp_02_21), .i_x4(w_pp_03_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_010), .ow_carry(w_c4to2_carry_23_010), .ow_cout(w_c4to2_cout_23_010)
);
wire w_c4to2_sum_23_011, w_c4to2_carry_23_011, w_c4to2_cout_23_011;
math_compressor_4to2 u_c4to2_23_011 (
    .i_x1(w_pp_04_19), .i_x2(w_pp_05_18),
    .i_x3(w_pp_06_17), .i_x4(w_pp_07_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_011), .ow_carry(w_c4to2_carry_23_011), .ow_cout(w_c4to2_cout_23_011)
);
wire w_c4to2_sum_23_012, w_c4to2_carry_23_012, w_c4to2_cout_23_012;
math_compressor_4to2 u_c4to2_23_012 (
    .i_x1(w_pp_08_15), .i_x2(w_pp_09_14),
    .i_x3(w_pp_10_13), .i_x4(w_pp_11_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_012), .ow_carry(w_c4to2_carry_23_012), .ow_cout(w_c4to2_cout_23_012)
);
wire w_c4to2_sum_23_013, w_c4to2_carry_23_013, w_c4to2_cout_23_013;
math_compressor_4to2 u_c4to2_23_013 (
    .i_x1(w_pp_12_11), .i_x2(w_pp_13_10),
    .i_x3(w_pp_14_09), .i_x4(w_pp_15_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_013), .ow_carry(w_c4to2_carry_23_013), .ow_cout(w_c4to2_cout_23_013)
);
wire w_c4to2_sum_23_014, w_c4to2_carry_23_014, w_c4to2_cout_23_014;
math_compressor_4to2 u_c4to2_23_014 (
    .i_x1(w_pp_16_07), .i_x2(w_pp_17_06),
    .i_x3(w_pp_18_05), .i_x4(w_pp_19_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_014), .ow_carry(w_c4to2_carry_23_014), .ow_cout(w_c4to2_cout_23_014)
);
wire w_c4to2_sum_24_015, w_c4to2_carry_24_015, w_c4to2_cout_24_015;
math_compressor_4to2 u_c4to2_24_015 (
    .i_x1(w_pp_01_23), .i_x2(w_pp_02_22),
    .i_x3(w_pp_03_21), .i_x4(w_pp_04_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_015), .ow_carry(w_c4to2_carry_24_015), .ow_cout(w_c4to2_cout_24_015)
);
wire w_c4to2_sum_24_016, w_c4to2_carry_24_016, w_c4to2_cout_24_016;
math_compressor_4to2 u_c4to2_24_016 (
    .i_x1(w_pp_05_19), .i_x2(w_pp_06_18),
    .i_x3(w_pp_07_17), .i_x4(w_pp_08_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_016), .ow_carry(w_c4to2_carry_24_016), .ow_cout(w_c4to2_cout_24_016)
);
wire w_c4to2_sum_24_017, w_c4to2_carry_24_017, w_c4to2_cout_24_017;
math_compressor_4to2 u_c4to2_24_017 (
    .i_x1(w_pp_09_15), .i_x2(w_pp_10_14),
    .i_x3(w_pp_11_13), .i_x4(w_pp_12_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_017), .ow_carry(w_c4to2_carry_24_017), .ow_cout(w_c4to2_cout_24_017)
);
wire w_c4to2_sum_24_018, w_c4to2_carry_24_018, w_c4to2_cout_24_018;
math_compressor_4to2 u_c4to2_24_018 (
    .i_x1(w_pp_13_11), .i_x2(w_pp_14_10),
    .i_x3(w_pp_15_09), .i_x4(w_pp_16_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_018), .ow_carry(w_c4to2_carry_24_018), .ow_cout(w_c4to2_cout_24_018)
);
wire w_c4to2_sum_24_019, w_c4to2_carry_24_019, w_c4to2_cout_24_019;
math_compressor_4to2 u_c4to2_24_019 (
    .i_x1(w_pp_17_07), .i_x2(w_pp_18_06),
    .i_x3(w_pp_19_05), .i_x4(w_pp_20_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_019), .ow_carry(w_c4to2_carry_24_019), .ow_cout(w_c4to2_cout_24_019)
);
wire w_c4to2_sum_25_020, w_c4to2_carry_25_020, w_c4to2_cout_25_020;
math_compressor_4to2 u_c4to2_25_020 (
    .i_x1(w_pp_02_23), .i_x2(w_pp_03_22),
    .i_x3(w_pp_04_21), .i_x4(w_pp_05_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_020), .ow_carry(w_c4to2_carry_25_020), .ow_cout(w_c4to2_cout_25_020)
);
wire w_c4to2_sum_25_021, w_c4to2_carry_25_021, w_c4to2_cout_25_021;
math_compressor_4to2 u_c4to2_25_021 (
    .i_x1(w_pp_06_19), .i_x2(w_pp_07_18),
    .i_x3(w_pp_08_17), .i_x4(w_pp_09_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_021), .ow_carry(w_c4to2_carry_25_021), .ow_cout(w_c4to2_cout_25_021)
);
wire w_c4to2_sum_25_022, w_c4to2_carry_25_022, w_c4to2_cout_25_022;
math_compressor_4to2 u_c4to2_25_022 (
    .i_x1(w_pp_10_15), .i_x2(w_pp_11_14),
    .i_x3(w_pp_12_13), .i_x4(w_pp_13_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_022), .ow_carry(w_c4to2_carry_25_022), .ow_cout(w_c4to2_cout_25_022)
);
wire w_c4to2_sum_25_023, w_c4to2_carry_25_023, w_c4to2_cout_25_023;
math_compressor_4to2 u_c4to2_25_023 (
    .i_x1(w_pp_14_11), .i_x2(w_pp_15_10),
    .i_x3(w_pp_16_09), .i_x4(w_pp_17_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_023), .ow_carry(w_c4to2_carry_25_023), .ow_cout(w_c4to2_cout_25_023)
);
wire w_c4to2_sum_25_024, w_c4to2_carry_25_024, w_c4to2_cout_25_024;
math_compressor_4to2 u_c4to2_25_024 (
    .i_x1(w_pp_18_07), .i_x2(w_pp_19_06),
    .i_x3(w_pp_20_05), .i_x4(w_pp_21_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_024), .ow_carry(w_c4to2_carry_25_024), .ow_cout(w_c4to2_cout_25_024)
);
wire w_c4to2_sum_26_025, w_c4to2_carry_26_025, w_c4to2_cout_26_025;
math_compressor_4to2 u_c4to2_26_025 (
    .i_x1(w_pp_03_23), .i_x2(w_pp_04_22),
    .i_x3(w_pp_05_21), .i_x4(w_pp_06_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_025), .ow_carry(w_c4to2_carry_26_025), .ow_cout(w_c4to2_cout_26_025)
);
wire w_c4to2_sum_26_026, w_c4to2_carry_26_026, w_c4to2_cout_26_026;
math_compressor_4to2 u_c4to2_26_026 (
    .i_x1(w_pp_07_19), .i_x2(w_pp_08_18),
    .i_x3(w_pp_09_17), .i_x4(w_pp_10_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_026), .ow_carry(w_c4to2_carry_26_026), .ow_cout(w_c4to2_cout_26_026)
);
wire w_c4to2_sum_26_027, w_c4to2_carry_26_027, w_c4to2_cout_26_027;
math_compressor_4to2 u_c4to2_26_027 (
    .i_x1(w_pp_11_15), .i_x2(w_pp_12_14),
    .i_x3(w_pp_13_13), .i_x4(w_pp_14_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_027), .ow_carry(w_c4to2_carry_26_027), .ow_cout(w_c4to2_cout_26_027)
);
wire w_c4to2_sum_26_028, w_c4to2_carry_26_028, w_c4to2_cout_26_028;
math_compressor_4to2 u_c4to2_26_028 (
    .i_x1(w_pp_15_11), .i_x2(w_pp_16_10),
    .i_x3(w_pp_17_09), .i_x4(w_pp_18_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_028), .ow_carry(w_c4to2_carry_26_028), .ow_cout(w_c4to2_cout_26_028)
);
wire w_c4to2_sum_27_029, w_c4to2_carry_27_029, w_c4to2_cout_27_029;
math_compressor_4to2 u_c4to2_27_029 (
    .i_x1(w_pp_04_23), .i_x2(w_pp_05_22),
    .i_x3(w_pp_06_21), .i_x4(w_pp_07_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_029), .ow_carry(w_c4to2_carry_27_029), .ow_cout(w_c4to2_cout_27_029)
);
wire w_c4to2_sum_27_030, w_c4to2_carry_27_030, w_c4to2_cout_27_030;
math_compressor_4to2 u_c4to2_27_030 (
    .i_x1(w_pp_08_19), .i_x2(w_pp_09_18),
    .i_x3(w_pp_10_17), .i_x4(w_pp_11_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_030), .ow_carry(w_c4to2_carry_27_030), .ow_cout(w_c4to2_cout_27_030)
);
wire w_c4to2_sum_27_031, w_c4to2_carry_27_031, w_c4to2_cout_27_031;
math_compressor_4to2 u_c4to2_27_031 (
    .i_x1(w_pp_12_15), .i_x2(w_pp_13_14),
    .i_x3(w_pp_14_13), .i_x4(w_pp_15_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_031), .ow_carry(w_c4to2_carry_27_031), .ow_cout(w_c4to2_cout_27_031)
);
wire w_c4to2_sum_28_032, w_c4to2_carry_28_032, w_c4to2_cout_28_032;
math_compressor_4to2 u_c4to2_28_032 (
    .i_x1(w_pp_05_23), .i_x2(w_pp_06_22),
    .i_x3(w_pp_07_21), .i_x4(w_pp_08_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_032), .ow_carry(w_c4to2_carry_28_032), .ow_cout(w_c4to2_cout_28_032)
);
wire w_c4to2_sum_28_033, w_c4to2_carry_28_033, w_c4to2_cout_28_033;
math_compressor_4to2 u_c4to2_28_033 (
    .i_x1(w_pp_09_19), .i_x2(w_pp_10_18),
    .i_x3(w_pp_11_17), .i_x4(w_pp_12_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_033), .ow_carry(w_c4to2_carry_28_033), .ow_cout(w_c4to2_cout_28_033)
);
wire w_c4to2_sum_29_034, w_c4to2_carry_29_034, w_c4to2_cout_29_034;
math_compressor_4to2 u_c4to2_29_034 (
    .i_x1(w_pp_06_23), .i_x2(w_pp_07_22),
    .i_x3(w_pp_08_21), .i_x4(w_pp_09_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_034), .ow_carry(w_c4to2_carry_29_034), .ow_cout(w_c4to2_cout_29_034)
);

// Dadda Reduction Stage 2: height 19 -> 13

wire w_c4to2_sum_13_035, w_c4to2_carry_13_035, w_c4to2_cout_13_035;
math_compressor_4to2 u_c4to2_13_035 (
    .i_x1(w_pp_00_13), .i_x2(w_pp_01_12),
    .i_x3(w_pp_02_11), .i_x4(w_pp_03_10),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_035), .ow_carry(w_c4to2_carry_13_035), .ow_cout(w_c4to2_cout_13_035)
);
wire w_c4to2_sum_14_036, w_c4to2_carry_14_036, w_c4to2_cout_14_036;
math_compressor_4to2 u_c4to2_14_036 (
    .i_x1(w_pp_00_14), .i_x2(w_pp_01_13),
    .i_x3(w_pp_02_12), .i_x4(w_pp_03_11),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_036), .ow_carry(w_c4to2_carry_14_036), .ow_cout(w_c4to2_cout_14_036)
);
wire w_c4to2_sum_14_037, w_c4to2_carry_14_037, w_c4to2_cout_14_037;
math_compressor_4to2 u_c4to2_14_037 (
    .i_x1(w_pp_04_10), .i_x2(w_pp_05_09),
    .i_x3(w_pp_06_08), .i_x4(w_pp_07_07),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_037), .ow_carry(w_c4to2_carry_14_037), .ow_cout(w_c4to2_cout_14_037)
);
wire w_c4to2_sum_15_038, w_c4to2_carry_15_038, w_c4to2_cout_15_038;
math_compressor_4to2 u_c4to2_15_038 (
    .i_x1(w_pp_00_15), .i_x2(w_pp_01_14),
    .i_x3(w_pp_02_13), .i_x4(w_pp_03_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_038), .ow_carry(w_c4to2_carry_15_038), .ow_cout(w_c4to2_cout_15_038)
);
wire w_c4to2_sum_15_039, w_c4to2_carry_15_039, w_c4to2_cout_15_039;
math_compressor_4to2 u_c4to2_15_039 (
    .i_x1(w_pp_04_11), .i_x2(w_pp_05_10),
    .i_x3(w_pp_06_09), .i_x4(w_pp_07_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_039), .ow_carry(w_c4to2_carry_15_039), .ow_cout(w_c4to2_cout_15_039)
);
wire w_c4to2_sum_15_040, w_c4to2_carry_15_040, w_c4to2_cout_15_040;
math_compressor_4to2 u_c4to2_15_040 (
    .i_x1(w_pp_08_07), .i_x2(w_pp_09_06),
    .i_x3(w_pp_10_05), .i_x4(w_pp_11_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_040), .ow_carry(w_c4to2_carry_15_040), .ow_cout(w_c4to2_cout_15_040)
);
wire w_c4to2_sum_16_041, w_c4to2_carry_16_041, w_c4to2_cout_16_041;
math_compressor_4to2 u_c4to2_16_041 (
    .i_x1(w_pp_00_16), .i_x2(w_pp_01_15),
    .i_x3(w_pp_02_14), .i_x4(w_pp_03_13),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_041), .ow_carry(w_c4to2_carry_16_041), .ow_cout(w_c4to2_cout_16_041)
);
wire w_c4to2_sum_16_042, w_c4to2_carry_16_042, w_c4to2_cout_16_042;
math_compressor_4to2 u_c4to2_16_042 (
    .i_x1(w_pp_04_12), .i_x2(w_pp_05_11),
    .i_x3(w_pp_06_10), .i_x4(w_pp_07_09),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_042), .ow_carry(w_c4to2_carry_16_042), .ow_cout(w_c4to2_cout_16_042)
);
wire w_c4to2_sum_16_043, w_c4to2_carry_16_043, w_c4to2_cout_16_043;
math_compressor_4to2 u_c4to2_16_043 (
    .i_x1(w_pp_08_08), .i_x2(w_pp_09_07),
    .i_x3(w_pp_10_06), .i_x4(w_pp_11_05),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_043), .ow_carry(w_c4to2_carry_16_043), .ow_cout(w_c4to2_cout_16_043)
);
wire w_c4to2_sum_16_044, w_c4to2_carry_16_044, w_c4to2_cout_16_044;
math_compressor_4to2 u_c4to2_16_044 (
    .i_x1(w_pp_12_04), .i_x2(w_pp_13_03),
    .i_x3(w_pp_14_02), .i_x4(w_pp_15_01),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_044), .ow_carry(w_c4to2_carry_16_044), .ow_cout(w_c4to2_cout_16_044)
);
wire w_c4to2_sum_17_045, w_c4to2_carry_17_045, w_c4to2_cout_17_045;
math_compressor_4to2 u_c4to2_17_045 (
    .i_x1(w_pp_00_17), .i_x2(w_pp_01_16),
    .i_x3(w_pp_02_15), .i_x4(w_pp_03_14),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_045), .ow_carry(w_c4to2_carry_17_045), .ow_cout(w_c4to2_cout_17_045)
);
wire w_c4to2_sum_17_046, w_c4to2_carry_17_046, w_c4to2_cout_17_046;
math_compressor_4to2 u_c4to2_17_046 (
    .i_x1(w_pp_04_13), .i_x2(w_pp_05_12),
    .i_x3(w_pp_06_11), .i_x4(w_pp_07_10),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_046), .ow_carry(w_c4to2_carry_17_046), .ow_cout(w_c4to2_cout_17_046)
);
wire w_c4to2_sum_17_047, w_c4to2_carry_17_047, w_c4to2_cout_17_047;
math_compressor_4to2 u_c4to2_17_047 (
    .i_x1(w_pp_08_09), .i_x2(w_pp_09_08),
    .i_x3(w_pp_10_07), .i_x4(w_pp_11_06),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_047), .ow_carry(w_c4to2_carry_17_047), .ow_cout(w_c4to2_cout_17_047)
);
wire w_c4to2_sum_17_048, w_c4to2_carry_17_048, w_c4to2_cout_17_048;
math_compressor_4to2 u_c4to2_17_048 (
    .i_x1(w_pp_12_05), .i_x2(w_pp_13_04),
    .i_x3(w_pp_14_03), .i_x4(w_pp_15_02),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_048), .ow_carry(w_c4to2_carry_17_048), .ow_cout(w_c4to2_cout_17_048)
);
wire w_c4to2_sum_17_049, w_c4to2_carry_17_049, w_c4to2_cout_17_049;
math_compressor_4to2 u_c4to2_17_049 (
    .i_x1(w_pp_16_01), .i_x2(w_pp_17_00),
    .i_x3(w_c4to2_carry_16_041), .i_x4(w_c4to2_cout_16_041),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_049), .ow_carry(w_c4to2_carry_17_049), .ow_cout(w_c4to2_cout_17_049)
);
wire w_c4to2_sum_18_050, w_c4to2_carry_18_050, w_c4to2_cout_18_050;
math_compressor_4to2 u_c4to2_18_050 (
    .i_x1(w_pp_00_18), .i_x2(w_pp_01_17),
    .i_x3(w_pp_02_16), .i_x4(w_pp_03_15),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_050), .ow_carry(w_c4to2_carry_18_050), .ow_cout(w_c4to2_cout_18_050)
);
wire w_c4to2_sum_18_051, w_c4to2_carry_18_051, w_c4to2_cout_18_051;
math_compressor_4to2 u_c4to2_18_051 (
    .i_x1(w_pp_04_14), .i_x2(w_pp_05_13),
    .i_x3(w_pp_06_12), .i_x4(w_pp_07_11),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_051), .ow_carry(w_c4to2_carry_18_051), .ow_cout(w_c4to2_cout_18_051)
);
wire w_c4to2_sum_18_052, w_c4to2_carry_18_052, w_c4to2_cout_18_052;
math_compressor_4to2 u_c4to2_18_052 (
    .i_x1(w_pp_08_10), .i_x2(w_pp_09_09),
    .i_x3(w_pp_10_08), .i_x4(w_pp_11_07),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_052), .ow_carry(w_c4to2_carry_18_052), .ow_cout(w_c4to2_cout_18_052)
);
wire w_c4to2_sum_18_053, w_c4to2_carry_18_053, w_c4to2_cout_18_053;
math_compressor_4to2 u_c4to2_18_053 (
    .i_x1(w_pp_12_06), .i_x2(w_pp_13_05),
    .i_x3(w_pp_14_04), .i_x4(w_pp_15_03),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_053), .ow_carry(w_c4to2_carry_18_053), .ow_cout(w_c4to2_cout_18_053)
);
wire w_c4to2_sum_18_054, w_c4to2_carry_18_054, w_c4to2_cout_18_054;
math_compressor_4to2 u_c4to2_18_054 (
    .i_x1(w_pp_16_02), .i_x2(w_pp_17_01),
    .i_x3(w_pp_18_00), .i_x4(w_c4to2_carry_17_045),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_054), .ow_carry(w_c4to2_carry_18_054), .ow_cout(w_c4to2_cout_18_054)
);
wire w_c4to2_sum_18_055, w_c4to2_carry_18_055, w_c4to2_cout_18_055;
math_compressor_4to2 u_c4to2_18_055 (
    .i_x1(w_c4to2_cout_17_045), .i_x2(w_c4to2_carry_17_046),
    .i_x3(w_c4to2_cout_17_046), .i_x4(w_c4to2_carry_17_047),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_055), .ow_carry(w_c4to2_carry_18_055), .ow_cout(w_c4to2_cout_18_055)
);
wire w_c4to2_sum_19_056, w_c4to2_carry_19_056, w_c4to2_cout_19_056;
math_compressor_4to2 u_c4to2_19_056 (
    .i_x1(w_pp_04_15), .i_x2(w_pp_05_14),
    .i_x3(w_pp_06_13), .i_x4(w_pp_07_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_056), .ow_carry(w_c4to2_carry_19_056), .ow_cout(w_c4to2_cout_19_056)
);
wire w_c4to2_sum_19_057, w_c4to2_carry_19_057, w_c4to2_cout_19_057;
math_compressor_4to2 u_c4to2_19_057 (
    .i_x1(w_pp_08_11), .i_x2(w_pp_09_10),
    .i_x3(w_pp_10_09), .i_x4(w_pp_11_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_057), .ow_carry(w_c4to2_carry_19_057), .ow_cout(w_c4to2_cout_19_057)
);
wire w_c4to2_sum_19_058, w_c4to2_carry_19_058, w_c4to2_cout_19_058;
math_compressor_4to2 u_c4to2_19_058 (
    .i_x1(w_pp_12_07), .i_x2(w_pp_13_06),
    .i_x3(w_pp_14_05), .i_x4(w_pp_15_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_058), .ow_carry(w_c4to2_carry_19_058), .ow_cout(w_c4to2_cout_19_058)
);
wire w_c4to2_sum_19_059, w_c4to2_carry_19_059, w_c4to2_cout_19_059;
math_compressor_4to2 u_c4to2_19_059 (
    .i_x1(w_pp_16_03), .i_x2(w_pp_17_02),
    .i_x3(w_pp_18_01), .i_x4(w_pp_19_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_059), .ow_carry(w_c4to2_carry_19_059), .ow_cout(w_c4to2_cout_19_059)
);
wire w_c4to2_sum_19_060, w_c4to2_carry_19_060, w_c4to2_cout_19_060;
math_compressor_4to2 u_c4to2_19_060 (
    .i_x1(w_c4to2_sum_19_000), .i_x2(w_c4to2_carry_18_050),
    .i_x3(w_c4to2_cout_18_050), .i_x4(w_c4to2_carry_18_051),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_060), .ow_carry(w_c4to2_carry_19_060), .ow_cout(w_c4to2_cout_19_060)
);
wire w_c4to2_sum_19_061, w_c4to2_carry_19_061, w_c4to2_cout_19_061;
math_compressor_4to2 u_c4to2_19_061 (
    .i_x1(w_c4to2_cout_18_051), .i_x2(w_c4to2_carry_18_052),
    .i_x3(w_c4to2_cout_18_052), .i_x4(w_c4to2_carry_18_053),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_061), .ow_carry(w_c4to2_carry_19_061), .ow_cout(w_c4to2_cout_19_061)
);
wire w_c4to2_sum_20_062, w_c4to2_carry_20_062, w_c4to2_cout_20_062;
math_compressor_4to2 u_c4to2_20_062 (
    .i_x1(w_pp_08_12), .i_x2(w_pp_09_11),
    .i_x3(w_pp_10_10), .i_x4(w_pp_11_09),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_062), .ow_carry(w_c4to2_carry_20_062), .ow_cout(w_c4to2_cout_20_062)
);
wire w_c4to2_sum_20_063, w_c4to2_carry_20_063, w_c4to2_cout_20_063;
math_compressor_4to2 u_c4to2_20_063 (
    .i_x1(w_pp_12_08), .i_x2(w_pp_13_07),
    .i_x3(w_pp_14_06), .i_x4(w_pp_15_05),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_063), .ow_carry(w_c4to2_carry_20_063), .ow_cout(w_c4to2_cout_20_063)
);
wire w_c4to2_sum_20_064, w_c4to2_carry_20_064, w_c4to2_cout_20_064;
math_compressor_4to2 u_c4to2_20_064 (
    .i_x1(w_pp_16_04), .i_x2(w_pp_17_03),
    .i_x3(w_pp_18_02), .i_x4(w_pp_19_01),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_064), .ow_carry(w_c4to2_carry_20_064), .ow_cout(w_c4to2_cout_20_064)
);
wire w_c4to2_sum_20_065, w_c4to2_carry_20_065, w_c4to2_cout_20_065;
math_compressor_4to2 u_c4to2_20_065 (
    .i_x1(w_pp_20_00), .i_x2(w_c4to2_carry_19_000),
    .i_x3(w_c4to2_cout_19_000), .i_x4(w_c4to2_sum_20_001),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_065), .ow_carry(w_c4to2_carry_20_065), .ow_cout(w_c4to2_cout_20_065)
);
wire w_c4to2_sum_20_066, w_c4to2_carry_20_066, w_c4to2_cout_20_066;
math_compressor_4to2 u_c4to2_20_066 (
    .i_x1(w_c4to2_sum_20_002), .i_x2(w_c4to2_carry_19_056),
    .i_x3(w_c4to2_cout_19_056), .i_x4(w_c4to2_carry_19_057),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_066), .ow_carry(w_c4to2_carry_20_066), .ow_cout(w_c4to2_cout_20_066)
);
wire w_c4to2_sum_20_067, w_c4to2_carry_20_067, w_c4to2_cout_20_067;
math_compressor_4to2 u_c4to2_20_067 (
    .i_x1(w_c4to2_cout_19_057), .i_x2(w_c4to2_carry_19_058),
    .i_x3(w_c4to2_cout_19_058), .i_x4(w_c4to2_carry_19_059),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_067), .ow_carry(w_c4to2_carry_20_067), .ow_cout(w_c4to2_cout_20_067)
);
wire w_c4to2_sum_21_068, w_c4to2_carry_21_068, w_c4to2_cout_21_068;
math_compressor_4to2 u_c4to2_21_068 (
    .i_x1(w_pp_12_09), .i_x2(w_pp_13_08),
    .i_x3(w_pp_14_07), .i_x4(w_pp_15_06),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_068), .ow_carry(w_c4to2_carry_21_068), .ow_cout(w_c4to2_cout_21_068)
);
wire w_c4to2_sum_21_069, w_c4to2_carry_21_069, w_c4to2_cout_21_069;
math_compressor_4to2 u_c4to2_21_069 (
    .i_x1(w_pp_16_05), .i_x2(w_pp_17_04),
    .i_x3(w_pp_18_03), .i_x4(w_pp_19_02),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_069), .ow_carry(w_c4to2_carry_21_069), .ow_cout(w_c4to2_cout_21_069)
);
wire w_c4to2_sum_21_070, w_c4to2_carry_21_070, w_c4to2_cout_21_070;
math_compressor_4to2 u_c4to2_21_070 (
    .i_x1(w_pp_20_01), .i_x2(w_pp_21_00),
    .i_x3(w_c4to2_carry_20_001), .i_x4(w_c4to2_cout_20_001),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_070), .ow_carry(w_c4to2_carry_21_070), .ow_cout(w_c4to2_cout_21_070)
);
wire w_c4to2_sum_21_071, w_c4to2_carry_21_071, w_c4to2_cout_21_071;
math_compressor_4to2 u_c4to2_21_071 (
    .i_x1(w_c4to2_carry_20_002), .i_x2(w_c4to2_cout_20_002),
    .i_x3(w_c4to2_sum_21_003), .i_x4(w_c4to2_sum_21_004),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_071), .ow_carry(w_c4to2_carry_21_071), .ow_cout(w_c4to2_cout_21_071)
);
wire w_c4to2_sum_21_072, w_c4to2_carry_21_072, w_c4to2_cout_21_072;
math_compressor_4to2 u_c4to2_21_072 (
    .i_x1(w_c4to2_sum_21_005), .i_x2(w_c4to2_carry_20_062),
    .i_x3(w_c4to2_cout_20_062), .i_x4(w_c4to2_carry_20_063),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_072), .ow_carry(w_c4to2_carry_21_072), .ow_cout(w_c4to2_cout_21_072)
);
wire w_c4to2_sum_21_073, w_c4to2_carry_21_073, w_c4to2_cout_21_073;
math_compressor_4to2 u_c4to2_21_073 (
    .i_x1(w_c4to2_cout_20_063), .i_x2(w_c4to2_carry_20_064),
    .i_x3(w_c4to2_cout_20_064), .i_x4(w_c4to2_carry_20_065),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_073), .ow_carry(w_c4to2_carry_21_073), .ow_cout(w_c4to2_cout_21_073)
);
wire w_c4to2_sum_22_074, w_c4to2_carry_22_074, w_c4to2_cout_22_074;
math_compressor_4to2 u_c4to2_22_074 (
    .i_x1(w_pp_16_06), .i_x2(w_pp_17_05),
    .i_x3(w_pp_18_04), .i_x4(w_pp_19_03),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_074), .ow_carry(w_c4to2_carry_22_074), .ow_cout(w_c4to2_cout_22_074)
);
wire w_c4to2_sum_22_075, w_c4to2_carry_22_075, w_c4to2_cout_22_075;
math_compressor_4to2 u_c4to2_22_075 (
    .i_x1(w_pp_20_02), .i_x2(w_pp_21_01),
    .i_x3(w_pp_22_00), .i_x4(w_c4to2_carry_21_003),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_075), .ow_carry(w_c4to2_carry_22_075), .ow_cout(w_c4to2_cout_22_075)
);
wire w_c4to2_sum_22_076, w_c4to2_carry_22_076, w_c4to2_cout_22_076;
math_compressor_4to2 u_c4to2_22_076 (
    .i_x1(w_c4to2_cout_21_003), .i_x2(w_c4to2_carry_21_004),
    .i_x3(w_c4to2_cout_21_004), .i_x4(w_c4to2_carry_21_005),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_076), .ow_carry(w_c4to2_carry_22_076), .ow_cout(w_c4to2_cout_22_076)
);
wire w_c4to2_sum_22_077, w_c4to2_carry_22_077, w_c4to2_cout_22_077;
math_compressor_4to2 u_c4to2_22_077 (
    .i_x1(w_c4to2_cout_21_005), .i_x2(w_c4to2_sum_22_006),
    .i_x3(w_c4to2_sum_22_007), .i_x4(w_c4to2_sum_22_008),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_077), .ow_carry(w_c4to2_carry_22_077), .ow_cout(w_c4to2_cout_22_077)
);
wire w_c4to2_sum_22_078, w_c4to2_carry_22_078, w_c4to2_cout_22_078;
math_compressor_4to2 u_c4to2_22_078 (
    .i_x1(w_c4to2_sum_22_009), .i_x2(w_c4to2_carry_21_068),
    .i_x3(w_c4to2_cout_21_068), .i_x4(w_c4to2_carry_21_069),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_078), .ow_carry(w_c4to2_carry_22_078), .ow_cout(w_c4to2_cout_22_078)
);
wire w_c4to2_sum_22_079, w_c4to2_carry_22_079, w_c4to2_cout_22_079;
math_compressor_4to2 u_c4to2_22_079 (
    .i_x1(w_c4to2_cout_21_069), .i_x2(w_c4to2_carry_21_070),
    .i_x3(w_c4to2_cout_21_070), .i_x4(w_c4to2_carry_21_071),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_079), .ow_carry(w_c4to2_carry_22_079), .ow_cout(w_c4to2_cout_22_079)
);
wire w_c4to2_sum_23_080, w_c4to2_carry_23_080, w_c4to2_cout_23_080;
math_compressor_4to2 u_c4to2_23_080 (
    .i_x1(w_pp_20_03), .i_x2(w_pp_21_02),
    .i_x3(w_pp_22_01), .i_x4(w_pp_23_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_080), .ow_carry(w_c4to2_carry_23_080), .ow_cout(w_c4to2_cout_23_080)
);
wire w_c4to2_sum_23_081, w_c4to2_carry_23_081, w_c4to2_cout_23_081;
math_compressor_4to2 u_c4to2_23_081 (
    .i_x1(w_c4to2_carry_22_006), .i_x2(w_c4to2_cout_22_006),
    .i_x3(w_c4to2_carry_22_007), .i_x4(w_c4to2_cout_22_007),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_081), .ow_carry(w_c4to2_carry_23_081), .ow_cout(w_c4to2_cout_23_081)
);
wire w_c4to2_sum_23_082, w_c4to2_carry_23_082, w_c4to2_cout_23_082;
math_compressor_4to2 u_c4to2_23_082 (
    .i_x1(w_c4to2_carry_22_008), .i_x2(w_c4to2_cout_22_008),
    .i_x3(w_c4to2_carry_22_009), .i_x4(w_c4to2_cout_22_009),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_082), .ow_carry(w_c4to2_carry_23_082), .ow_cout(w_c4to2_cout_23_082)
);
wire w_c4to2_sum_23_083, w_c4to2_carry_23_083, w_c4to2_cout_23_083;
math_compressor_4to2 u_c4to2_23_083 (
    .i_x1(w_c4to2_sum_23_010), .i_x2(w_c4to2_sum_23_011),
    .i_x3(w_c4to2_sum_23_012), .i_x4(w_c4to2_sum_23_013),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_083), .ow_carry(w_c4to2_carry_23_083), .ow_cout(w_c4to2_cout_23_083)
);
wire w_c4to2_sum_23_084, w_c4to2_carry_23_084, w_c4to2_cout_23_084;
math_compressor_4to2 u_c4to2_23_084 (
    .i_x1(w_c4to2_sum_23_014), .i_x2(w_c4to2_carry_22_074),
    .i_x3(w_c4to2_cout_22_074), .i_x4(w_c4to2_carry_22_075),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_084), .ow_carry(w_c4to2_carry_23_084), .ow_cout(w_c4to2_cout_23_084)
);
wire w_c4to2_sum_23_085, w_c4to2_carry_23_085, w_c4to2_cout_23_085;
math_compressor_4to2 u_c4to2_23_085 (
    .i_x1(w_c4to2_cout_22_075), .i_x2(w_c4to2_carry_22_076),
    .i_x3(w_c4to2_cout_22_076), .i_x4(w_c4to2_carry_22_077),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_085), .ow_carry(w_c4to2_carry_23_085), .ow_cout(w_c4to2_cout_23_085)
);
wire w_c4to2_sum_24_086, w_c4to2_carry_24_086, w_c4to2_cout_24_086;
math_compressor_4to2 u_c4to2_24_086 (
    .i_x1(w_pp_21_03), .i_x2(w_pp_22_02),
    .i_x3(w_pp_23_01), .i_x4(w_c4to2_carry_23_010),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_086), .ow_carry(w_c4to2_carry_24_086), .ow_cout(w_c4to2_cout_24_086)
);
wire w_c4to2_sum_24_087, w_c4to2_carry_24_087, w_c4to2_cout_24_087;
math_compressor_4to2 u_c4to2_24_087 (
    .i_x1(w_c4to2_cout_23_010), .i_x2(w_c4to2_carry_23_011),
    .i_x3(w_c4to2_cout_23_011), .i_x4(w_c4to2_carry_23_012),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_087), .ow_carry(w_c4to2_carry_24_087), .ow_cout(w_c4to2_cout_24_087)
);
wire w_c4to2_sum_24_088, w_c4to2_carry_24_088, w_c4to2_cout_24_088;
math_compressor_4to2 u_c4to2_24_088 (
    .i_x1(w_c4to2_cout_23_012), .i_x2(w_c4to2_carry_23_013),
    .i_x3(w_c4to2_cout_23_013), .i_x4(w_c4to2_carry_23_014),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_088), .ow_carry(w_c4to2_carry_24_088), .ow_cout(w_c4to2_cout_24_088)
);
wire w_c4to2_sum_24_089, w_c4to2_carry_24_089, w_c4to2_cout_24_089;
math_compressor_4to2 u_c4to2_24_089 (
    .i_x1(w_c4to2_cout_23_014), .i_x2(w_c4to2_sum_24_015),
    .i_x3(w_c4to2_sum_24_016), .i_x4(w_c4to2_sum_24_017),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_089), .ow_carry(w_c4to2_carry_24_089), .ow_cout(w_c4to2_cout_24_089)
);
wire w_c4to2_sum_24_090, w_c4to2_carry_24_090, w_c4to2_cout_24_090;
math_compressor_4to2 u_c4to2_24_090 (
    .i_x1(w_c4to2_sum_24_018), .i_x2(w_c4to2_sum_24_019),
    .i_x3(w_c4to2_carry_23_080), .i_x4(w_c4to2_cout_23_080),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_090), .ow_carry(w_c4to2_carry_24_090), .ow_cout(w_c4to2_cout_24_090)
);
wire w_c4to2_sum_24_091, w_c4to2_carry_24_091, w_c4to2_cout_24_091;
math_compressor_4to2 u_c4to2_24_091 (
    .i_x1(w_c4to2_carry_23_081), .i_x2(w_c4to2_cout_23_081),
    .i_x3(w_c4to2_carry_23_082), .i_x4(w_c4to2_cout_23_082),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_091), .ow_carry(w_c4to2_carry_24_091), .ow_cout(w_c4to2_cout_24_091)
);
wire w_c4to2_sum_25_092, w_c4to2_carry_25_092, w_c4to2_cout_25_092;
math_compressor_4to2 u_c4to2_25_092 (
    .i_x1(w_pp_22_03), .i_x2(w_pp_23_02),
    .i_x3(w_c4to2_carry_24_015), .i_x4(w_c4to2_cout_24_015),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_092), .ow_carry(w_c4to2_carry_25_092), .ow_cout(w_c4to2_cout_25_092)
);
wire w_c4to2_sum_25_093, w_c4to2_carry_25_093, w_c4to2_cout_25_093;
math_compressor_4to2 u_c4to2_25_093 (
    .i_x1(w_c4to2_carry_24_016), .i_x2(w_c4to2_cout_24_016),
    .i_x3(w_c4to2_carry_24_017), .i_x4(w_c4to2_cout_24_017),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_093), .ow_carry(w_c4to2_carry_25_093), .ow_cout(w_c4to2_cout_25_093)
);
wire w_c4to2_sum_25_094, w_c4to2_carry_25_094, w_c4to2_cout_25_094;
math_compressor_4to2 u_c4to2_25_094 (
    .i_x1(w_c4to2_carry_24_018), .i_x2(w_c4to2_cout_24_018),
    .i_x3(w_c4to2_carry_24_019), .i_x4(w_c4to2_cout_24_019),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_094), .ow_carry(w_c4to2_carry_25_094), .ow_cout(w_c4to2_cout_25_094)
);
wire w_c4to2_sum_25_095, w_c4to2_carry_25_095, w_c4to2_cout_25_095;
math_compressor_4to2 u_c4to2_25_095 (
    .i_x1(w_c4to2_sum_25_020), .i_x2(w_c4to2_sum_25_021),
    .i_x3(w_c4to2_sum_25_022), .i_x4(w_c4to2_sum_25_023),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_095), .ow_carry(w_c4to2_carry_25_095), .ow_cout(w_c4to2_cout_25_095)
);
wire w_c4to2_sum_25_096, w_c4to2_carry_25_096, w_c4to2_cout_25_096;
math_compressor_4to2 u_c4to2_25_096 (
    .i_x1(w_c4to2_sum_25_024), .i_x2(w_c4to2_carry_24_086),
    .i_x3(w_c4to2_cout_24_086), .i_x4(w_c4to2_carry_24_087),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_096), .ow_carry(w_c4to2_carry_25_096), .ow_cout(w_c4to2_cout_25_096)
);
wire w_c4to2_sum_25_097, w_c4to2_carry_25_097, w_c4to2_cout_25_097;
math_compressor_4to2 u_c4to2_25_097 (
    .i_x1(w_c4to2_cout_24_087), .i_x2(w_c4to2_carry_24_088),
    .i_x3(w_c4to2_cout_24_088), .i_x4(w_c4to2_carry_24_089),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_097), .ow_carry(w_c4to2_carry_25_097), .ow_cout(w_c4to2_cout_25_097)
);
wire w_c4to2_sum_26_098, w_c4to2_carry_26_098, w_c4to2_cout_26_098;
math_compressor_4to2 u_c4to2_26_098 (
    .i_x1(w_pp_19_07), .i_x2(w_pp_20_06),
    .i_x3(w_pp_21_05), .i_x4(w_pp_22_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_098), .ow_carry(w_c4to2_carry_26_098), .ow_cout(w_c4to2_cout_26_098)
);
wire w_c4to2_sum_26_099, w_c4to2_carry_26_099, w_c4to2_cout_26_099;
math_compressor_4to2 u_c4to2_26_099 (
    .i_x1(w_pp_23_03), .i_x2(w_c4to2_carry_25_020),
    .i_x3(w_c4to2_cout_25_020), .i_x4(w_c4to2_carry_25_021),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_099), .ow_carry(w_c4to2_carry_26_099), .ow_cout(w_c4to2_cout_26_099)
);
wire w_c4to2_sum_26_100, w_c4to2_carry_26_100, w_c4to2_cout_26_100;
math_compressor_4to2 u_c4to2_26_100 (
    .i_x1(w_c4to2_cout_25_021), .i_x2(w_c4to2_carry_25_022),
    .i_x3(w_c4to2_cout_25_022), .i_x4(w_c4to2_carry_25_023),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_100), .ow_carry(w_c4to2_carry_26_100), .ow_cout(w_c4to2_cout_26_100)
);
wire w_c4to2_sum_26_101, w_c4to2_carry_26_101, w_c4to2_cout_26_101;
math_compressor_4to2 u_c4to2_26_101 (
    .i_x1(w_c4to2_cout_25_023), .i_x2(w_c4to2_carry_25_024),
    .i_x3(w_c4to2_cout_25_024), .i_x4(w_c4to2_sum_26_025),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_101), .ow_carry(w_c4to2_carry_26_101), .ow_cout(w_c4to2_cout_26_101)
);
wire w_c4to2_sum_26_102, w_c4to2_carry_26_102, w_c4to2_cout_26_102;
math_compressor_4to2 u_c4to2_26_102 (
    .i_x1(w_c4to2_sum_26_026), .i_x2(w_c4to2_sum_26_027),
    .i_x3(w_c4to2_sum_26_028), .i_x4(w_c4to2_carry_25_092),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_102), .ow_carry(w_c4to2_carry_26_102), .ow_cout(w_c4to2_cout_26_102)
);
wire w_c4to2_sum_26_103, w_c4to2_carry_26_103, w_c4to2_cout_26_103;
math_compressor_4to2 u_c4to2_26_103 (
    .i_x1(w_c4to2_cout_25_092), .i_x2(w_c4to2_carry_25_093),
    .i_x3(w_c4to2_cout_25_093), .i_x4(w_c4to2_carry_25_094),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_103), .ow_carry(w_c4to2_carry_26_103), .ow_cout(w_c4to2_cout_26_103)
);
wire w_c4to2_sum_27_104, w_c4to2_carry_27_104, w_c4to2_cout_27_104;
math_compressor_4to2 u_c4to2_27_104 (
    .i_x1(w_pp_16_11), .i_x2(w_pp_17_10),
    .i_x3(w_pp_18_09), .i_x4(w_pp_19_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_104), .ow_carry(w_c4to2_carry_27_104), .ow_cout(w_c4to2_cout_27_104)
);
wire w_c4to2_sum_27_105, w_c4to2_carry_27_105, w_c4to2_cout_27_105;
math_compressor_4to2 u_c4to2_27_105 (
    .i_x1(w_pp_20_07), .i_x2(w_pp_21_06),
    .i_x3(w_pp_22_05), .i_x4(w_pp_23_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_105), .ow_carry(w_c4to2_carry_27_105), .ow_cout(w_c4to2_cout_27_105)
);
wire w_c4to2_sum_27_106, w_c4to2_carry_27_106, w_c4to2_cout_27_106;
math_compressor_4to2 u_c4to2_27_106 (
    .i_x1(w_c4to2_carry_26_025), .i_x2(w_c4to2_cout_26_025),
    .i_x3(w_c4to2_carry_26_026), .i_x4(w_c4to2_cout_26_026),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_106), .ow_carry(w_c4to2_carry_27_106), .ow_cout(w_c4to2_cout_27_106)
);
wire w_c4to2_sum_27_107, w_c4to2_carry_27_107, w_c4to2_cout_27_107;
math_compressor_4to2 u_c4to2_27_107 (
    .i_x1(w_c4to2_carry_26_027), .i_x2(w_c4to2_cout_26_027),
    .i_x3(w_c4to2_carry_26_028), .i_x4(w_c4to2_cout_26_028),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_107), .ow_carry(w_c4to2_carry_27_107), .ow_cout(w_c4to2_cout_27_107)
);
wire w_c4to2_sum_27_108, w_c4to2_carry_27_108, w_c4to2_cout_27_108;
math_compressor_4to2 u_c4to2_27_108 (
    .i_x1(w_c4to2_sum_27_029), .i_x2(w_c4to2_sum_27_030),
    .i_x3(w_c4to2_sum_27_031), .i_x4(w_c4to2_carry_26_098),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_108), .ow_carry(w_c4to2_carry_27_108), .ow_cout(w_c4to2_cout_27_108)
);
wire w_c4to2_sum_27_109, w_c4to2_carry_27_109, w_c4to2_cout_27_109;
math_compressor_4to2 u_c4to2_27_109 (
    .i_x1(w_c4to2_cout_26_098), .i_x2(w_c4to2_carry_26_099),
    .i_x3(w_c4to2_cout_26_099), .i_x4(w_c4to2_carry_26_100),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_109), .ow_carry(w_c4to2_carry_27_109), .ow_cout(w_c4to2_cout_27_109)
);
wire w_c4to2_sum_28_110, w_c4to2_carry_28_110, w_c4to2_cout_28_110;
math_compressor_4to2 u_c4to2_28_110 (
    .i_x1(w_pp_13_15), .i_x2(w_pp_14_14),
    .i_x3(w_pp_15_13), .i_x4(w_pp_16_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_110), .ow_carry(w_c4to2_carry_28_110), .ow_cout(w_c4to2_cout_28_110)
);
wire w_c4to2_sum_28_111, w_c4to2_carry_28_111, w_c4to2_cout_28_111;
math_compressor_4to2 u_c4to2_28_111 (
    .i_x1(w_pp_17_11), .i_x2(w_pp_18_10),
    .i_x3(w_pp_19_09), .i_x4(w_pp_20_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_111), .ow_carry(w_c4to2_carry_28_111), .ow_cout(w_c4to2_cout_28_111)
);
wire w_c4to2_sum_28_112, w_c4to2_carry_28_112, w_c4to2_cout_28_112;
math_compressor_4to2 u_c4to2_28_112 (
    .i_x1(w_pp_21_07), .i_x2(w_pp_22_06),
    .i_x3(w_pp_23_05), .i_x4(w_c4to2_carry_27_029),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_112), .ow_carry(w_c4to2_carry_28_112), .ow_cout(w_c4to2_cout_28_112)
);
wire w_c4to2_sum_28_113, w_c4to2_carry_28_113, w_c4to2_cout_28_113;
math_compressor_4to2 u_c4to2_28_113 (
    .i_x1(w_c4to2_cout_27_029), .i_x2(w_c4to2_carry_27_030),
    .i_x3(w_c4to2_cout_27_030), .i_x4(w_c4to2_carry_27_031),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_113), .ow_carry(w_c4to2_carry_28_113), .ow_cout(w_c4to2_cout_28_113)
);
wire w_c4to2_sum_28_114, w_c4to2_carry_28_114, w_c4to2_cout_28_114;
math_compressor_4to2 u_c4to2_28_114 (
    .i_x1(w_c4to2_cout_27_031), .i_x2(w_c4to2_sum_28_032),
    .i_x3(w_c4to2_sum_28_033), .i_x4(w_c4to2_carry_27_104),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_114), .ow_carry(w_c4to2_carry_28_114), .ow_cout(w_c4to2_cout_28_114)
);
wire w_c4to2_sum_28_115, w_c4to2_carry_28_115, w_c4to2_cout_28_115;
math_compressor_4to2 u_c4to2_28_115 (
    .i_x1(w_c4to2_cout_27_104), .i_x2(w_c4to2_carry_27_105),
    .i_x3(w_c4to2_cout_27_105), .i_x4(w_c4to2_carry_27_106),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_115), .ow_carry(w_c4to2_carry_28_115), .ow_cout(w_c4to2_cout_28_115)
);
wire w_c4to2_sum_29_116, w_c4to2_carry_29_116, w_c4to2_cout_29_116;
math_compressor_4to2 u_c4to2_29_116 (
    .i_x1(w_pp_10_19), .i_x2(w_pp_11_18),
    .i_x3(w_pp_12_17), .i_x4(w_pp_13_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_116), .ow_carry(w_c4to2_carry_29_116), .ow_cout(w_c4to2_cout_29_116)
);
wire w_c4to2_sum_29_117, w_c4to2_carry_29_117, w_c4to2_cout_29_117;
math_compressor_4to2 u_c4to2_29_117 (
    .i_x1(w_pp_14_15), .i_x2(w_pp_15_14),
    .i_x3(w_pp_16_13), .i_x4(w_pp_17_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_117), .ow_carry(w_c4to2_carry_29_117), .ow_cout(w_c4to2_cout_29_117)
);
wire w_c4to2_sum_29_118, w_c4to2_carry_29_118, w_c4to2_cout_29_118;
math_compressor_4to2 u_c4to2_29_118 (
    .i_x1(w_pp_18_11), .i_x2(w_pp_19_10),
    .i_x3(w_pp_20_09), .i_x4(w_pp_21_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_118), .ow_carry(w_c4to2_carry_29_118), .ow_cout(w_c4to2_cout_29_118)
);
wire w_c4to2_sum_29_119, w_c4to2_carry_29_119, w_c4to2_cout_29_119;
math_compressor_4to2 u_c4to2_29_119 (
    .i_x1(w_pp_22_07), .i_x2(w_pp_23_06),
    .i_x3(w_c4to2_carry_28_032), .i_x4(w_c4to2_cout_28_032),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_119), .ow_carry(w_c4to2_carry_29_119), .ow_cout(w_c4to2_cout_29_119)
);
wire w_c4to2_sum_29_120, w_c4to2_carry_29_120, w_c4to2_cout_29_120;
math_compressor_4to2 u_c4to2_29_120 (
    .i_x1(w_c4to2_carry_28_033), .i_x2(w_c4to2_cout_28_033),
    .i_x3(w_c4to2_sum_29_034), .i_x4(w_c4to2_carry_28_110),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_120), .ow_carry(w_c4to2_carry_29_120), .ow_cout(w_c4to2_cout_29_120)
);
wire w_c4to2_sum_29_121, w_c4to2_carry_29_121, w_c4to2_cout_29_121;
math_compressor_4to2 u_c4to2_29_121 (
    .i_x1(w_c4to2_cout_28_110), .i_x2(w_c4to2_carry_28_111),
    .i_x3(w_c4to2_cout_28_111), .i_x4(w_c4to2_carry_28_112),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_121), .ow_carry(w_c4to2_carry_29_121), .ow_cout(w_c4to2_cout_29_121)
);
wire w_c4to2_sum_30_122, w_c4to2_carry_30_122, w_c4to2_cout_30_122;
math_compressor_4to2 u_c4to2_30_122 (
    .i_x1(w_pp_07_23), .i_x2(w_pp_08_22),
    .i_x3(w_pp_09_21), .i_x4(w_pp_10_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_122), .ow_carry(w_c4to2_carry_30_122), .ow_cout(w_c4to2_cout_30_122)
);
wire w_c4to2_sum_30_123, w_c4to2_carry_30_123, w_c4to2_cout_30_123;
math_compressor_4to2 u_c4to2_30_123 (
    .i_x1(w_pp_11_19), .i_x2(w_pp_12_18),
    .i_x3(w_pp_13_17), .i_x4(w_pp_14_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_123), .ow_carry(w_c4to2_carry_30_123), .ow_cout(w_c4to2_cout_30_123)
);
wire w_c4to2_sum_30_124, w_c4to2_carry_30_124, w_c4to2_cout_30_124;
math_compressor_4to2 u_c4to2_30_124 (
    .i_x1(w_pp_15_15), .i_x2(w_pp_16_14),
    .i_x3(w_pp_17_13), .i_x4(w_pp_18_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_124), .ow_carry(w_c4to2_carry_30_124), .ow_cout(w_c4to2_cout_30_124)
);
wire w_c4to2_sum_30_125, w_c4to2_carry_30_125, w_c4to2_cout_30_125;
math_compressor_4to2 u_c4to2_30_125 (
    .i_x1(w_pp_19_11), .i_x2(w_pp_20_10),
    .i_x3(w_pp_21_09), .i_x4(w_pp_22_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_125), .ow_carry(w_c4to2_carry_30_125), .ow_cout(w_c4to2_cout_30_125)
);
wire w_c4to2_sum_30_126, w_c4to2_carry_30_126, w_c4to2_cout_30_126;
math_compressor_4to2 u_c4to2_30_126 (
    .i_x1(w_pp_23_07), .i_x2(w_c4to2_carry_29_034),
    .i_x3(w_c4to2_cout_29_034), .i_x4(w_c4to2_carry_29_116),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_126), .ow_carry(w_c4to2_carry_30_126), .ow_cout(w_c4to2_cout_30_126)
);
wire w_c4to2_sum_30_127, w_c4to2_carry_30_127, w_c4to2_cout_30_127;
math_compressor_4to2 u_c4to2_30_127 (
    .i_x1(w_c4to2_cout_29_116), .i_x2(w_c4to2_carry_29_117),
    .i_x3(w_c4to2_cout_29_117), .i_x4(w_c4to2_carry_29_118),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_127), .ow_carry(w_c4to2_carry_30_127), .ow_cout(w_c4to2_cout_30_127)
);
wire w_c4to2_sum_31_128, w_c4to2_carry_31_128, w_c4to2_cout_31_128;
math_compressor_4to2 u_c4to2_31_128 (
    .i_x1(w_pp_08_23), .i_x2(w_pp_09_22),
    .i_x3(w_pp_10_21), .i_x4(w_pp_11_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_128), .ow_carry(w_c4to2_carry_31_128), .ow_cout(w_c4to2_cout_31_128)
);
wire w_c4to2_sum_31_129, w_c4to2_carry_31_129, w_c4to2_cout_31_129;
math_compressor_4to2 u_c4to2_31_129 (
    .i_x1(w_pp_12_19), .i_x2(w_pp_13_18),
    .i_x3(w_pp_14_17), .i_x4(w_pp_15_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_129), .ow_carry(w_c4to2_carry_31_129), .ow_cout(w_c4to2_cout_31_129)
);
wire w_c4to2_sum_31_130, w_c4to2_carry_31_130, w_c4to2_cout_31_130;
math_compressor_4to2 u_c4to2_31_130 (
    .i_x1(w_pp_16_15), .i_x2(w_pp_17_14),
    .i_x3(w_pp_18_13), .i_x4(w_pp_19_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_130), .ow_carry(w_c4to2_carry_31_130), .ow_cout(w_c4to2_cout_31_130)
);
wire w_c4to2_sum_31_131, w_c4to2_carry_31_131, w_c4to2_cout_31_131;
math_compressor_4to2 u_c4to2_31_131 (
    .i_x1(w_pp_20_11), .i_x2(w_pp_21_10),
    .i_x3(w_pp_22_09), .i_x4(w_pp_23_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_131), .ow_carry(w_c4to2_carry_31_131), .ow_cout(w_c4to2_cout_31_131)
);
wire w_c4to2_sum_31_132, w_c4to2_carry_31_132, w_c4to2_cout_31_132;
math_compressor_4to2 u_c4to2_31_132 (
    .i_x1(w_c4to2_carry_30_122), .i_x2(w_c4to2_cout_30_122),
    .i_x3(w_c4to2_carry_30_123), .i_x4(w_c4to2_cout_30_123),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_132), .ow_carry(w_c4to2_carry_31_132), .ow_cout(w_c4to2_cout_31_132)
);
wire w_c4to2_sum_32_133, w_c4to2_carry_32_133, w_c4to2_cout_32_133;
math_compressor_4to2 u_c4to2_32_133 (
    .i_x1(w_pp_09_23), .i_x2(w_pp_10_22),
    .i_x3(w_pp_11_21), .i_x4(w_pp_12_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_133), .ow_carry(w_c4to2_carry_32_133), .ow_cout(w_c4to2_cout_32_133)
);
wire w_c4to2_sum_32_134, w_c4to2_carry_32_134, w_c4to2_cout_32_134;
math_compressor_4to2 u_c4to2_32_134 (
    .i_x1(w_pp_13_19), .i_x2(w_pp_14_18),
    .i_x3(w_pp_15_17), .i_x4(w_pp_16_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_134), .ow_carry(w_c4to2_carry_32_134), .ow_cout(w_c4to2_cout_32_134)
);
wire w_c4to2_sum_32_135, w_c4to2_carry_32_135, w_c4to2_cout_32_135;
math_compressor_4to2 u_c4to2_32_135 (
    .i_x1(w_pp_17_15), .i_x2(w_pp_18_14),
    .i_x3(w_pp_19_13), .i_x4(w_pp_20_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_135), .ow_carry(w_c4to2_carry_32_135), .ow_cout(w_c4to2_cout_32_135)
);
wire w_c4to2_sum_32_136, w_c4to2_carry_32_136, w_c4to2_cout_32_136;
math_compressor_4to2 u_c4to2_32_136 (
    .i_x1(w_pp_21_11), .i_x2(w_pp_22_10),
    .i_x3(w_pp_23_09), .i_x4(w_c4to2_carry_31_128),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_136), .ow_carry(w_c4to2_carry_32_136), .ow_cout(w_c4to2_cout_32_136)
);
wire w_c4to2_sum_33_137, w_c4to2_carry_33_137, w_c4to2_cout_33_137;
math_compressor_4to2 u_c4to2_33_137 (
    .i_x1(w_pp_10_23), .i_x2(w_pp_11_22),
    .i_x3(w_pp_12_21), .i_x4(w_pp_13_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_137), .ow_carry(w_c4to2_carry_33_137), .ow_cout(w_c4to2_cout_33_137)
);
wire w_c4to2_sum_33_138, w_c4to2_carry_33_138, w_c4to2_cout_33_138;
math_compressor_4to2 u_c4to2_33_138 (
    .i_x1(w_pp_14_19), .i_x2(w_pp_15_18),
    .i_x3(w_pp_16_17), .i_x4(w_pp_17_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_138), .ow_carry(w_c4to2_carry_33_138), .ow_cout(w_c4to2_cout_33_138)
);
wire w_c4to2_sum_33_139, w_c4to2_carry_33_139, w_c4to2_cout_33_139;
math_compressor_4to2 u_c4to2_33_139 (
    .i_x1(w_pp_18_15), .i_x2(w_pp_19_14),
    .i_x3(w_pp_20_13), .i_x4(w_pp_21_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_139), .ow_carry(w_c4to2_carry_33_139), .ow_cout(w_c4to2_cout_33_139)
);
wire w_c4to2_sum_34_140, w_c4to2_carry_34_140, w_c4to2_cout_34_140;
math_compressor_4to2 u_c4to2_34_140 (
    .i_x1(w_pp_11_23), .i_x2(w_pp_12_22),
    .i_x3(w_pp_13_21), .i_x4(w_pp_14_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_140), .ow_carry(w_c4to2_carry_34_140), .ow_cout(w_c4to2_cout_34_140)
);
wire w_c4to2_sum_34_141, w_c4to2_carry_34_141, w_c4to2_cout_34_141;
math_compressor_4to2 u_c4to2_34_141 (
    .i_x1(w_pp_15_19), .i_x2(w_pp_16_18),
    .i_x3(w_pp_17_17), .i_x4(w_pp_18_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_141), .ow_carry(w_c4to2_carry_34_141), .ow_cout(w_c4to2_cout_34_141)
);
wire w_c4to2_sum_35_142, w_c4to2_carry_35_142, w_c4to2_cout_35_142;
math_compressor_4to2 u_c4to2_35_142 (
    .i_x1(w_pp_12_23), .i_x2(w_pp_13_22),
    .i_x3(w_pp_14_21), .i_x4(w_pp_15_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_142), .ow_carry(w_c4to2_carry_35_142), .ow_cout(w_c4to2_cout_35_142)
);

// Dadda Reduction Stage 3: height 13 -> 9

wire w_c4to2_sum_09_143, w_c4to2_carry_09_143, w_c4to2_cout_09_143;
math_compressor_4to2 u_c4to2_09_143 (
    .i_x1(w_pp_00_09), .i_x2(w_pp_01_08),
    .i_x3(w_pp_02_07), .i_x4(w_pp_03_06),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_143), .ow_carry(w_c4to2_carry_09_143), .ow_cout(w_c4to2_cout_09_143)
);
wire w_c4to2_sum_10_144, w_c4to2_carry_10_144, w_c4to2_cout_10_144;
math_compressor_4to2 u_c4to2_10_144 (
    .i_x1(w_pp_00_10), .i_x2(w_pp_01_09),
    .i_x3(w_pp_02_08), .i_x4(w_pp_03_07),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_144), .ow_carry(w_c4to2_carry_10_144), .ow_cout(w_c4to2_cout_10_144)
);
wire w_c4to2_sum_10_145, w_c4to2_carry_10_145, w_c4to2_cout_10_145;
math_compressor_4to2 u_c4to2_10_145 (
    .i_x1(w_pp_04_06), .i_x2(w_pp_05_05),
    .i_x3(w_pp_06_04), .i_x4(w_pp_07_03),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_145), .ow_carry(w_c4to2_carry_10_145), .ow_cout(w_c4to2_cout_10_145)
);
wire w_c4to2_sum_11_146, w_c4to2_carry_11_146, w_c4to2_cout_11_146;
math_compressor_4to2 u_c4to2_11_146 (
    .i_x1(w_pp_00_11), .i_x2(w_pp_01_10),
    .i_x3(w_pp_02_09), .i_x4(w_pp_03_08),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_146), .ow_carry(w_c4to2_carry_11_146), .ow_cout(w_c4to2_cout_11_146)
);
wire w_c4to2_sum_11_147, w_c4to2_carry_11_147, w_c4to2_cout_11_147;
math_compressor_4to2 u_c4to2_11_147 (
    .i_x1(w_pp_04_07), .i_x2(w_pp_05_06),
    .i_x3(w_pp_06_05), .i_x4(w_pp_07_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_147), .ow_carry(w_c4to2_carry_11_147), .ow_cout(w_c4to2_cout_11_147)
);
wire w_c4to2_sum_11_148, w_c4to2_carry_11_148, w_c4to2_cout_11_148;
math_compressor_4to2 u_c4to2_11_148 (
    .i_x1(w_pp_08_03), .i_x2(w_pp_09_02),
    .i_x3(w_pp_10_01), .i_x4(w_pp_11_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_148), .ow_carry(w_c4to2_carry_11_148), .ow_cout(w_c4to2_cout_11_148)
);
wire w_c4to2_sum_12_149, w_c4to2_carry_12_149, w_c4to2_cout_12_149;
math_compressor_4to2 u_c4to2_12_149 (
    .i_x1(w_pp_00_12), .i_x2(w_pp_01_11),
    .i_x3(w_pp_02_10), .i_x4(w_pp_03_09),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_149), .ow_carry(w_c4to2_carry_12_149), .ow_cout(w_c4to2_cout_12_149)
);
wire w_c4to2_sum_12_150, w_c4to2_carry_12_150, w_c4to2_cout_12_150;
math_compressor_4to2 u_c4to2_12_150 (
    .i_x1(w_pp_04_08), .i_x2(w_pp_05_07),
    .i_x3(w_pp_06_06), .i_x4(w_pp_07_05),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_150), .ow_carry(w_c4to2_carry_12_150), .ow_cout(w_c4to2_cout_12_150)
);
wire w_c4to2_sum_12_151, w_c4to2_carry_12_151, w_c4to2_cout_12_151;
math_compressor_4to2 u_c4to2_12_151 (
    .i_x1(w_pp_08_04), .i_x2(w_pp_09_03),
    .i_x3(w_pp_10_02), .i_x4(w_pp_11_01),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_151), .ow_carry(w_c4to2_carry_12_151), .ow_cout(w_c4to2_cout_12_151)
);
wire w_c4to2_sum_12_152, w_c4to2_carry_12_152, w_c4to2_cout_12_152;
math_compressor_4to2 u_c4to2_12_152 (
    .i_x1(w_pp_12_00), .i_x2(w_c4to2_carry_11_146),
    .i_x3(w_c4to2_cout_11_146), .i_x4(w_c4to2_carry_11_147),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_152), .ow_carry(w_c4to2_carry_12_152), .ow_cout(w_c4to2_cout_12_152)
);
wire w_c4to2_sum_13_153, w_c4to2_carry_13_153, w_c4to2_cout_13_153;
math_compressor_4to2 u_c4to2_13_153 (
    .i_x1(w_pp_04_09), .i_x2(w_pp_05_08),
    .i_x3(w_pp_06_07), .i_x4(w_pp_07_06),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_153), .ow_carry(w_c4to2_carry_13_153), .ow_cout(w_c4to2_cout_13_153)
);
wire w_c4to2_sum_13_154, w_c4to2_carry_13_154, w_c4to2_cout_13_154;
math_compressor_4to2 u_c4to2_13_154 (
    .i_x1(w_pp_08_05), .i_x2(w_pp_09_04),
    .i_x3(w_pp_10_03), .i_x4(w_pp_11_02),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_154), .ow_carry(w_c4to2_carry_13_154), .ow_cout(w_c4to2_cout_13_154)
);
wire w_c4to2_sum_13_155, w_c4to2_carry_13_155, w_c4to2_cout_13_155;
math_compressor_4to2 u_c4to2_13_155 (
    .i_x1(w_pp_12_01), .i_x2(w_pp_13_00),
    .i_x3(w_c4to2_sum_13_035), .i_x4(w_c4to2_carry_12_149),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_155), .ow_carry(w_c4to2_carry_13_155), .ow_cout(w_c4to2_cout_13_155)
);
wire w_c4to2_sum_13_156, w_c4to2_carry_13_156, w_c4to2_cout_13_156;
math_compressor_4to2 u_c4to2_13_156 (
    .i_x1(w_c4to2_cout_12_149), .i_x2(w_c4to2_carry_12_150),
    .i_x3(w_c4to2_cout_12_150), .i_x4(w_c4to2_carry_12_151),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_156), .ow_carry(w_c4to2_carry_13_156), .ow_cout(w_c4to2_cout_13_156)
);
wire w_c4to2_sum_14_157, w_c4to2_carry_14_157, w_c4to2_cout_14_157;
math_compressor_4to2 u_c4to2_14_157 (
    .i_x1(w_pp_08_06), .i_x2(w_pp_09_05),
    .i_x3(w_pp_10_04), .i_x4(w_pp_11_03),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_157), .ow_carry(w_c4to2_carry_14_157), .ow_cout(w_c4to2_cout_14_157)
);
wire w_c4to2_sum_14_158, w_c4to2_carry_14_158, w_c4to2_cout_14_158;
math_compressor_4to2 u_c4to2_14_158 (
    .i_x1(w_pp_12_02), .i_x2(w_pp_13_01),
    .i_x3(w_pp_14_00), .i_x4(w_c4to2_carry_13_035),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_158), .ow_carry(w_c4to2_carry_14_158), .ow_cout(w_c4to2_cout_14_158)
);
wire w_c4to2_sum_14_159, w_c4to2_carry_14_159, w_c4to2_cout_14_159;
math_compressor_4to2 u_c4to2_14_159 (
    .i_x1(w_c4to2_cout_13_035), .i_x2(w_c4to2_sum_14_036),
    .i_x3(w_c4to2_sum_14_037), .i_x4(w_c4to2_carry_13_153),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_159), .ow_carry(w_c4to2_carry_14_159), .ow_cout(w_c4to2_cout_14_159)
);
wire w_c4to2_sum_14_160, w_c4to2_carry_14_160, w_c4to2_cout_14_160;
math_compressor_4to2 u_c4to2_14_160 (
    .i_x1(w_c4to2_cout_13_153), .i_x2(w_c4to2_carry_13_154),
    .i_x3(w_c4to2_cout_13_154), .i_x4(w_c4to2_carry_13_155),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_160), .ow_carry(w_c4to2_carry_14_160), .ow_cout(w_c4to2_cout_14_160)
);
wire w_c4to2_sum_15_161, w_c4to2_carry_15_161, w_c4to2_cout_15_161;
math_compressor_4to2 u_c4to2_15_161 (
    .i_x1(w_pp_12_03), .i_x2(w_pp_13_02),
    .i_x3(w_pp_14_01), .i_x4(w_pp_15_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_161), .ow_carry(w_c4to2_carry_15_161), .ow_cout(w_c4to2_cout_15_161)
);
wire w_c4to2_sum_15_162, w_c4to2_carry_15_162, w_c4to2_cout_15_162;
math_compressor_4to2 u_c4to2_15_162 (
    .i_x1(w_c4to2_carry_14_036), .i_x2(w_c4to2_cout_14_036),
    .i_x3(w_c4to2_carry_14_037), .i_x4(w_c4to2_cout_14_037),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_162), .ow_carry(w_c4to2_carry_15_162), .ow_cout(w_c4to2_cout_15_162)
);
wire w_c4to2_sum_15_163, w_c4to2_carry_15_163, w_c4to2_cout_15_163;
math_compressor_4to2 u_c4to2_15_163 (
    .i_x1(w_c4to2_sum_15_038), .i_x2(w_c4to2_sum_15_039),
    .i_x3(w_c4to2_sum_15_040), .i_x4(w_c4to2_carry_14_157),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_163), .ow_carry(w_c4to2_carry_15_163), .ow_cout(w_c4to2_cout_15_163)
);
wire w_c4to2_sum_15_164, w_c4to2_carry_15_164, w_c4to2_cout_15_164;
math_compressor_4to2 u_c4to2_15_164 (
    .i_x1(w_c4to2_cout_14_157), .i_x2(w_c4to2_carry_14_158),
    .i_x3(w_c4to2_cout_14_158), .i_x4(w_c4to2_carry_14_159),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_164), .ow_carry(w_c4to2_carry_15_164), .ow_cout(w_c4to2_cout_15_164)
);
wire w_c4to2_sum_16_165, w_c4to2_carry_16_165, w_c4to2_cout_16_165;
math_compressor_4to2 u_c4to2_16_165 (
    .i_x1(w_pp_16_00), .i_x2(w_c4to2_carry_15_038),
    .i_x3(w_c4to2_cout_15_038), .i_x4(w_c4to2_carry_15_039),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_165), .ow_carry(w_c4to2_carry_16_165), .ow_cout(w_c4to2_cout_16_165)
);
wire w_c4to2_sum_16_166, w_c4to2_carry_16_166, w_c4to2_cout_16_166;
math_compressor_4to2 u_c4to2_16_166 (
    .i_x1(w_c4to2_cout_15_039), .i_x2(w_c4to2_carry_15_040),
    .i_x3(w_c4to2_cout_15_040), .i_x4(w_c4to2_sum_16_041),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_166), .ow_carry(w_c4to2_carry_16_166), .ow_cout(w_c4to2_cout_16_166)
);
wire w_c4to2_sum_16_167, w_c4to2_carry_16_167, w_c4to2_cout_16_167;
math_compressor_4to2 u_c4to2_16_167 (
    .i_x1(w_c4to2_sum_16_042), .i_x2(w_c4to2_sum_16_043),
    .i_x3(w_c4to2_sum_16_044), .i_x4(w_c4to2_carry_15_161),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_167), .ow_carry(w_c4to2_carry_16_167), .ow_cout(w_c4to2_cout_16_167)
);
wire w_c4to2_sum_16_168, w_c4to2_carry_16_168, w_c4to2_cout_16_168;
math_compressor_4to2 u_c4to2_16_168 (
    .i_x1(w_c4to2_cout_15_161), .i_x2(w_c4to2_carry_15_162),
    .i_x3(w_c4to2_cout_15_162), .i_x4(w_c4to2_carry_15_163),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_168), .ow_carry(w_c4to2_carry_16_168), .ow_cout(w_c4to2_cout_16_168)
);
wire w_c4to2_sum_17_169, w_c4to2_carry_17_169, w_c4to2_cout_17_169;
math_compressor_4to2 u_c4to2_17_169 (
    .i_x1(w_c4to2_carry_16_042), .i_x2(w_c4to2_cout_16_042),
    .i_x3(w_c4to2_carry_16_043), .i_x4(w_c4to2_cout_16_043),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_169), .ow_carry(w_c4to2_carry_17_169), .ow_cout(w_c4to2_cout_17_169)
);
wire w_c4to2_sum_17_170, w_c4to2_carry_17_170, w_c4to2_cout_17_170;
math_compressor_4to2 u_c4to2_17_170 (
    .i_x1(w_c4to2_carry_16_044), .i_x2(w_c4to2_cout_16_044),
    .i_x3(w_c4to2_sum_17_045), .i_x4(w_c4to2_sum_17_046),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_170), .ow_carry(w_c4to2_carry_17_170), .ow_cout(w_c4to2_cout_17_170)
);
wire w_c4to2_sum_17_171, w_c4to2_carry_17_171, w_c4to2_cout_17_171;
math_compressor_4to2 u_c4to2_17_171 (
    .i_x1(w_c4to2_sum_17_047), .i_x2(w_c4to2_sum_17_048),
    .i_x3(w_c4to2_sum_17_049), .i_x4(w_c4to2_carry_16_165),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_171), .ow_carry(w_c4to2_carry_17_171), .ow_cout(w_c4to2_cout_17_171)
);
wire w_c4to2_sum_17_172, w_c4to2_carry_17_172, w_c4to2_cout_17_172;
math_compressor_4to2 u_c4to2_17_172 (
    .i_x1(w_c4to2_cout_16_165), .i_x2(w_c4to2_carry_16_166),
    .i_x3(w_c4to2_cout_16_166), .i_x4(w_c4to2_carry_16_167),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_172), .ow_carry(w_c4to2_carry_17_172), .ow_cout(w_c4to2_cout_17_172)
);
wire w_c4to2_sum_18_173, w_c4to2_carry_18_173, w_c4to2_cout_18_173;
math_compressor_4to2 u_c4to2_18_173 (
    .i_x1(w_c4to2_cout_17_047), .i_x2(w_c4to2_carry_17_048),
    .i_x3(w_c4to2_cout_17_048), .i_x4(w_c4to2_carry_17_049),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_173), .ow_carry(w_c4to2_carry_18_173), .ow_cout(w_c4to2_cout_18_173)
);
wire w_c4to2_sum_18_174, w_c4to2_carry_18_174, w_c4to2_cout_18_174;
math_compressor_4to2 u_c4to2_18_174 (
    .i_x1(w_c4to2_cout_17_049), .i_x2(w_c4to2_sum_18_050),
    .i_x3(w_c4to2_sum_18_051), .i_x4(w_c4to2_sum_18_052),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_174), .ow_carry(w_c4to2_carry_18_174), .ow_cout(w_c4to2_cout_18_174)
);
wire w_c4to2_sum_18_175, w_c4to2_carry_18_175, w_c4to2_cout_18_175;
math_compressor_4to2 u_c4to2_18_175 (
    .i_x1(w_c4to2_sum_18_053), .i_x2(w_c4to2_sum_18_054),
    .i_x3(w_c4to2_sum_18_055), .i_x4(w_c4to2_carry_17_169),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_175), .ow_carry(w_c4to2_carry_18_175), .ow_cout(w_c4to2_cout_18_175)
);
wire w_c4to2_sum_18_176, w_c4to2_carry_18_176, w_c4to2_cout_18_176;
math_compressor_4to2 u_c4to2_18_176 (
    .i_x1(w_c4to2_cout_17_169), .i_x2(w_c4to2_carry_17_170),
    .i_x3(w_c4to2_cout_17_170), .i_x4(w_c4to2_carry_17_171),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_176), .ow_carry(w_c4to2_carry_18_176), .ow_cout(w_c4to2_cout_18_176)
);
wire w_c4to2_sum_19_177, w_c4to2_carry_19_177, w_c4to2_cout_19_177;
math_compressor_4to2 u_c4to2_19_177 (
    .i_x1(w_c4to2_cout_18_053), .i_x2(w_c4to2_carry_18_054),
    .i_x3(w_c4to2_cout_18_054), .i_x4(w_c4to2_carry_18_055),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_177), .ow_carry(w_c4to2_carry_19_177), .ow_cout(w_c4to2_cout_19_177)
);
wire w_c4to2_sum_19_178, w_c4to2_carry_19_178, w_c4to2_cout_19_178;
math_compressor_4to2 u_c4to2_19_178 (
    .i_x1(w_c4to2_cout_18_055), .i_x2(w_c4to2_sum_19_056),
    .i_x3(w_c4to2_sum_19_057), .i_x4(w_c4to2_sum_19_058),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_178), .ow_carry(w_c4to2_carry_19_178), .ow_cout(w_c4to2_cout_19_178)
);
wire w_c4to2_sum_19_179, w_c4to2_carry_19_179, w_c4to2_cout_19_179;
math_compressor_4to2 u_c4to2_19_179 (
    .i_x1(w_c4to2_sum_19_059), .i_x2(w_c4to2_sum_19_060),
    .i_x3(w_c4to2_sum_19_061), .i_x4(w_c4to2_carry_18_173),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_179), .ow_carry(w_c4to2_carry_19_179), .ow_cout(w_c4to2_cout_19_179)
);
wire w_c4to2_sum_19_180, w_c4to2_carry_19_180, w_c4to2_cout_19_180;
math_compressor_4to2 u_c4to2_19_180 (
    .i_x1(w_c4to2_cout_18_173), .i_x2(w_c4to2_carry_18_174),
    .i_x3(w_c4to2_cout_18_174), .i_x4(w_c4to2_carry_18_175),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_180), .ow_carry(w_c4to2_carry_19_180), .ow_cout(w_c4to2_cout_19_180)
);
wire w_c4to2_sum_20_181, w_c4to2_carry_20_181, w_c4to2_cout_20_181;
math_compressor_4to2 u_c4to2_20_181 (
    .i_x1(w_c4to2_cout_19_059), .i_x2(w_c4to2_carry_19_060),
    .i_x3(w_c4to2_cout_19_060), .i_x4(w_c4to2_carry_19_061),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_181), .ow_carry(w_c4to2_carry_20_181), .ow_cout(w_c4to2_cout_20_181)
);
wire w_c4to2_sum_20_182, w_c4to2_carry_20_182, w_c4to2_cout_20_182;
math_compressor_4to2 u_c4to2_20_182 (
    .i_x1(w_c4to2_cout_19_061), .i_x2(w_c4to2_sum_20_062),
    .i_x3(w_c4to2_sum_20_063), .i_x4(w_c4to2_sum_20_064),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_182), .ow_carry(w_c4to2_carry_20_182), .ow_cout(w_c4to2_cout_20_182)
);
wire w_c4to2_sum_20_183, w_c4to2_carry_20_183, w_c4to2_cout_20_183;
math_compressor_4to2 u_c4to2_20_183 (
    .i_x1(w_c4to2_sum_20_065), .i_x2(w_c4to2_sum_20_066),
    .i_x3(w_c4to2_sum_20_067), .i_x4(w_c4to2_carry_19_177),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_183), .ow_carry(w_c4to2_carry_20_183), .ow_cout(w_c4to2_cout_20_183)
);
wire w_c4to2_sum_20_184, w_c4to2_carry_20_184, w_c4to2_cout_20_184;
math_compressor_4to2 u_c4to2_20_184 (
    .i_x1(w_c4to2_cout_19_177), .i_x2(w_c4to2_carry_19_178),
    .i_x3(w_c4to2_cout_19_178), .i_x4(w_c4to2_carry_19_179),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_184), .ow_carry(w_c4to2_carry_20_184), .ow_cout(w_c4to2_cout_20_184)
);
wire w_c4to2_sum_21_185, w_c4to2_carry_21_185, w_c4to2_cout_21_185;
math_compressor_4to2 u_c4to2_21_185 (
    .i_x1(w_c4to2_cout_20_065), .i_x2(w_c4to2_carry_20_066),
    .i_x3(w_c4to2_cout_20_066), .i_x4(w_c4to2_carry_20_067),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_185), .ow_carry(w_c4to2_carry_21_185), .ow_cout(w_c4to2_cout_21_185)
);
wire w_c4to2_sum_21_186, w_c4to2_carry_21_186, w_c4to2_cout_21_186;
math_compressor_4to2 u_c4to2_21_186 (
    .i_x1(w_c4to2_cout_20_067), .i_x2(w_c4to2_sum_21_068),
    .i_x3(w_c4to2_sum_21_069), .i_x4(w_c4to2_sum_21_070),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_186), .ow_carry(w_c4to2_carry_21_186), .ow_cout(w_c4to2_cout_21_186)
);
wire w_c4to2_sum_21_187, w_c4to2_carry_21_187, w_c4to2_cout_21_187;
math_compressor_4to2 u_c4to2_21_187 (
    .i_x1(w_c4to2_sum_21_071), .i_x2(w_c4to2_sum_21_072),
    .i_x3(w_c4to2_sum_21_073), .i_x4(w_c4to2_carry_20_181),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_187), .ow_carry(w_c4to2_carry_21_187), .ow_cout(w_c4to2_cout_21_187)
);
wire w_c4to2_sum_21_188, w_c4to2_carry_21_188, w_c4to2_cout_21_188;
math_compressor_4to2 u_c4to2_21_188 (
    .i_x1(w_c4to2_cout_20_181), .i_x2(w_c4to2_carry_20_182),
    .i_x3(w_c4to2_cout_20_182), .i_x4(w_c4to2_carry_20_183),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_188), .ow_carry(w_c4to2_carry_21_188), .ow_cout(w_c4to2_cout_21_188)
);
wire w_c4to2_sum_22_189, w_c4to2_carry_22_189, w_c4to2_cout_22_189;
math_compressor_4to2 u_c4to2_22_189 (
    .i_x1(w_c4to2_cout_21_071), .i_x2(w_c4to2_carry_21_072),
    .i_x3(w_c4to2_cout_21_072), .i_x4(w_c4to2_carry_21_073),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_189), .ow_carry(w_c4to2_carry_22_189), .ow_cout(w_c4to2_cout_22_189)
);
wire w_c4to2_sum_22_190, w_c4to2_carry_22_190, w_c4to2_cout_22_190;
math_compressor_4to2 u_c4to2_22_190 (
    .i_x1(w_c4to2_cout_21_073), .i_x2(w_c4to2_sum_22_074),
    .i_x3(w_c4to2_sum_22_075), .i_x4(w_c4to2_sum_22_076),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_190), .ow_carry(w_c4to2_carry_22_190), .ow_cout(w_c4to2_cout_22_190)
);
wire w_c4to2_sum_22_191, w_c4to2_carry_22_191, w_c4to2_cout_22_191;
math_compressor_4to2 u_c4to2_22_191 (
    .i_x1(w_c4to2_sum_22_077), .i_x2(w_c4to2_sum_22_078),
    .i_x3(w_c4to2_sum_22_079), .i_x4(w_c4to2_carry_21_185),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_191), .ow_carry(w_c4to2_carry_22_191), .ow_cout(w_c4to2_cout_22_191)
);
wire w_c4to2_sum_22_192, w_c4to2_carry_22_192, w_c4to2_cout_22_192;
math_compressor_4to2 u_c4to2_22_192 (
    .i_x1(w_c4to2_cout_21_185), .i_x2(w_c4to2_carry_21_186),
    .i_x3(w_c4to2_cout_21_186), .i_x4(w_c4to2_carry_21_187),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_192), .ow_carry(w_c4to2_carry_22_192), .ow_cout(w_c4to2_cout_22_192)
);
wire w_c4to2_sum_23_193, w_c4to2_carry_23_193, w_c4to2_cout_23_193;
math_compressor_4to2 u_c4to2_23_193 (
    .i_x1(w_c4to2_cout_22_077), .i_x2(w_c4to2_carry_22_078),
    .i_x3(w_c4to2_cout_22_078), .i_x4(w_c4to2_carry_22_079),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_193), .ow_carry(w_c4to2_carry_23_193), .ow_cout(w_c4to2_cout_23_193)
);
wire w_c4to2_sum_23_194, w_c4to2_carry_23_194, w_c4to2_cout_23_194;
math_compressor_4to2 u_c4to2_23_194 (
    .i_x1(w_c4to2_cout_22_079), .i_x2(w_c4to2_sum_23_080),
    .i_x3(w_c4to2_sum_23_081), .i_x4(w_c4to2_sum_23_082),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_194), .ow_carry(w_c4to2_carry_23_194), .ow_cout(w_c4to2_cout_23_194)
);
wire w_c4to2_sum_23_195, w_c4to2_carry_23_195, w_c4to2_cout_23_195;
math_compressor_4to2 u_c4to2_23_195 (
    .i_x1(w_c4to2_sum_23_083), .i_x2(w_c4to2_sum_23_084),
    .i_x3(w_c4to2_sum_23_085), .i_x4(w_c4to2_carry_22_189),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_195), .ow_carry(w_c4to2_carry_23_195), .ow_cout(w_c4to2_cout_23_195)
);
wire w_c4to2_sum_23_196, w_c4to2_carry_23_196, w_c4to2_cout_23_196;
math_compressor_4to2 u_c4to2_23_196 (
    .i_x1(w_c4to2_cout_22_189), .i_x2(w_c4to2_carry_22_190),
    .i_x3(w_c4to2_cout_22_190), .i_x4(w_c4to2_carry_22_191),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_196), .ow_carry(w_c4to2_carry_23_196), .ow_cout(w_c4to2_cout_23_196)
);
wire w_c4to2_sum_24_197, w_c4to2_carry_24_197, w_c4to2_cout_24_197;
math_compressor_4to2 u_c4to2_24_197 (
    .i_x1(w_c4to2_carry_23_083), .i_x2(w_c4to2_cout_23_083),
    .i_x3(w_c4to2_carry_23_084), .i_x4(w_c4to2_cout_23_084),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_197), .ow_carry(w_c4to2_carry_24_197), .ow_cout(w_c4to2_cout_24_197)
);
wire w_c4to2_sum_24_198, w_c4to2_carry_24_198, w_c4to2_cout_24_198;
math_compressor_4to2 u_c4to2_24_198 (
    .i_x1(w_c4to2_carry_23_085), .i_x2(w_c4to2_cout_23_085),
    .i_x3(w_c4to2_sum_24_086), .i_x4(w_c4to2_sum_24_087),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_198), .ow_carry(w_c4to2_carry_24_198), .ow_cout(w_c4to2_cout_24_198)
);
wire w_c4to2_sum_24_199, w_c4to2_carry_24_199, w_c4to2_cout_24_199;
math_compressor_4to2 u_c4to2_24_199 (
    .i_x1(w_c4to2_sum_24_088), .i_x2(w_c4to2_sum_24_089),
    .i_x3(w_c4to2_sum_24_090), .i_x4(w_c4to2_sum_24_091),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_199), .ow_carry(w_c4to2_carry_24_199), .ow_cout(w_c4to2_cout_24_199)
);
wire w_c4to2_sum_24_200, w_c4to2_carry_24_200, w_c4to2_cout_24_200;
math_compressor_4to2 u_c4to2_24_200 (
    .i_x1(w_c4to2_carry_23_193), .i_x2(w_c4to2_cout_23_193),
    .i_x3(w_c4to2_carry_23_194), .i_x4(w_c4to2_cout_23_194),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_200), .ow_carry(w_c4to2_carry_24_200), .ow_cout(w_c4to2_cout_24_200)
);
wire w_c4to2_sum_25_201, w_c4to2_carry_25_201, w_c4to2_cout_25_201;
math_compressor_4to2 u_c4to2_25_201 (
    .i_x1(w_c4to2_cout_24_089), .i_x2(w_c4to2_carry_24_090),
    .i_x3(w_c4to2_cout_24_090), .i_x4(w_c4to2_carry_24_091),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_201), .ow_carry(w_c4to2_carry_25_201), .ow_cout(w_c4to2_cout_25_201)
);
wire w_c4to2_sum_25_202, w_c4to2_carry_25_202, w_c4to2_cout_25_202;
math_compressor_4to2 u_c4to2_25_202 (
    .i_x1(w_c4to2_cout_24_091), .i_x2(w_c4to2_sum_25_092),
    .i_x3(w_c4to2_sum_25_093), .i_x4(w_c4to2_sum_25_094),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_202), .ow_carry(w_c4to2_carry_25_202), .ow_cout(w_c4to2_cout_25_202)
);
wire w_c4to2_sum_25_203, w_c4to2_carry_25_203, w_c4to2_cout_25_203;
math_compressor_4to2 u_c4to2_25_203 (
    .i_x1(w_c4to2_sum_25_095), .i_x2(w_c4to2_sum_25_096),
    .i_x3(w_c4to2_sum_25_097), .i_x4(w_c4to2_carry_24_197),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_203), .ow_carry(w_c4to2_carry_25_203), .ow_cout(w_c4to2_cout_25_203)
);
wire w_c4to2_sum_25_204, w_c4to2_carry_25_204, w_c4to2_cout_25_204;
math_compressor_4to2 u_c4to2_25_204 (
    .i_x1(w_c4to2_cout_24_197), .i_x2(w_c4to2_carry_24_198),
    .i_x3(w_c4to2_cout_24_198), .i_x4(w_c4to2_carry_24_199),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_204), .ow_carry(w_c4to2_carry_25_204), .ow_cout(w_c4to2_cout_25_204)
);
wire w_c4to2_sum_26_205, w_c4to2_carry_26_205, w_c4to2_cout_26_205;
math_compressor_4to2 u_c4to2_26_205 (
    .i_x1(w_c4to2_cout_25_094), .i_x2(w_c4to2_carry_25_095),
    .i_x3(w_c4to2_cout_25_095), .i_x4(w_c4to2_carry_25_096),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_205), .ow_carry(w_c4to2_carry_26_205), .ow_cout(w_c4to2_cout_26_205)
);
wire w_c4to2_sum_26_206, w_c4to2_carry_26_206, w_c4to2_cout_26_206;
math_compressor_4to2 u_c4to2_26_206 (
    .i_x1(w_c4to2_cout_25_096), .i_x2(w_c4to2_carry_25_097),
    .i_x3(w_c4to2_cout_25_097), .i_x4(w_c4to2_sum_26_098),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_206), .ow_carry(w_c4to2_carry_26_206), .ow_cout(w_c4to2_cout_26_206)
);
wire w_c4to2_sum_26_207, w_c4to2_carry_26_207, w_c4to2_cout_26_207;
math_compressor_4to2 u_c4to2_26_207 (
    .i_x1(w_c4to2_sum_26_099), .i_x2(w_c4to2_sum_26_100),
    .i_x3(w_c4to2_sum_26_101), .i_x4(w_c4to2_sum_26_102),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_207), .ow_carry(w_c4to2_carry_26_207), .ow_cout(w_c4to2_cout_26_207)
);
wire w_c4to2_sum_26_208, w_c4to2_carry_26_208, w_c4to2_cout_26_208;
math_compressor_4to2 u_c4to2_26_208 (
    .i_x1(w_c4to2_sum_26_103), .i_x2(w_c4to2_carry_25_201),
    .i_x3(w_c4to2_cout_25_201), .i_x4(w_c4to2_carry_25_202),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_208), .ow_carry(w_c4to2_carry_26_208), .ow_cout(w_c4to2_cout_26_208)
);
wire w_c4to2_sum_27_209, w_c4to2_carry_27_209, w_c4to2_cout_27_209;
math_compressor_4to2 u_c4to2_27_209 (
    .i_x1(w_c4to2_cout_26_100), .i_x2(w_c4to2_carry_26_101),
    .i_x3(w_c4to2_cout_26_101), .i_x4(w_c4to2_carry_26_102),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_209), .ow_carry(w_c4to2_carry_27_209), .ow_cout(w_c4to2_cout_27_209)
);
wire w_c4to2_sum_27_210, w_c4to2_carry_27_210, w_c4to2_cout_27_210;
math_compressor_4to2 u_c4to2_27_210 (
    .i_x1(w_c4to2_cout_26_102), .i_x2(w_c4to2_carry_26_103),
    .i_x3(w_c4to2_cout_26_103), .i_x4(w_c4to2_sum_27_104),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_210), .ow_carry(w_c4to2_carry_27_210), .ow_cout(w_c4to2_cout_27_210)
);
wire w_c4to2_sum_27_211, w_c4to2_carry_27_211, w_c4to2_cout_27_211;
math_compressor_4to2 u_c4to2_27_211 (
    .i_x1(w_c4to2_sum_27_105), .i_x2(w_c4to2_sum_27_106),
    .i_x3(w_c4to2_sum_27_107), .i_x4(w_c4to2_sum_27_108),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_211), .ow_carry(w_c4to2_carry_27_211), .ow_cout(w_c4to2_cout_27_211)
);
wire w_c4to2_sum_27_212, w_c4to2_carry_27_212, w_c4to2_cout_27_212;
math_compressor_4to2 u_c4to2_27_212 (
    .i_x1(w_c4to2_sum_27_109), .i_x2(w_c4to2_carry_26_205),
    .i_x3(w_c4to2_cout_26_205), .i_x4(w_c4to2_carry_26_206),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_212), .ow_carry(w_c4to2_carry_27_212), .ow_cout(w_c4to2_cout_27_212)
);
wire w_c4to2_sum_28_213, w_c4to2_carry_28_213, w_c4to2_cout_28_213;
math_compressor_4to2 u_c4to2_28_213 (
    .i_x1(w_c4to2_cout_27_106), .i_x2(w_c4to2_carry_27_107),
    .i_x3(w_c4to2_cout_27_107), .i_x4(w_c4to2_carry_27_108),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_213), .ow_carry(w_c4to2_carry_28_213), .ow_cout(w_c4to2_cout_28_213)
);
wire w_c4to2_sum_28_214, w_c4to2_carry_28_214, w_c4to2_cout_28_214;
math_compressor_4to2 u_c4to2_28_214 (
    .i_x1(w_c4to2_cout_27_108), .i_x2(w_c4to2_carry_27_109),
    .i_x3(w_c4to2_cout_27_109), .i_x4(w_c4to2_sum_28_110),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_214), .ow_carry(w_c4to2_carry_28_214), .ow_cout(w_c4to2_cout_28_214)
);
wire w_c4to2_sum_28_215, w_c4to2_carry_28_215, w_c4to2_cout_28_215;
math_compressor_4to2 u_c4to2_28_215 (
    .i_x1(w_c4to2_sum_28_111), .i_x2(w_c4to2_sum_28_112),
    .i_x3(w_c4to2_sum_28_113), .i_x4(w_c4to2_sum_28_114),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_215), .ow_carry(w_c4to2_carry_28_215), .ow_cout(w_c4to2_cout_28_215)
);
wire w_c4to2_sum_28_216, w_c4to2_carry_28_216, w_c4to2_cout_28_216;
math_compressor_4to2 u_c4to2_28_216 (
    .i_x1(w_c4to2_sum_28_115), .i_x2(w_c4to2_carry_27_209),
    .i_x3(w_c4to2_cout_27_209), .i_x4(w_c4to2_carry_27_210),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_216), .ow_carry(w_c4to2_carry_28_216), .ow_cout(w_c4to2_cout_28_216)
);
wire w_c4to2_sum_29_217, w_c4to2_carry_29_217, w_c4to2_cout_29_217;
math_compressor_4to2 u_c4to2_29_217 (
    .i_x1(w_c4to2_cout_28_112), .i_x2(w_c4to2_carry_28_113),
    .i_x3(w_c4to2_cout_28_113), .i_x4(w_c4to2_carry_28_114),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_217), .ow_carry(w_c4to2_carry_29_217), .ow_cout(w_c4to2_cout_29_217)
);
wire w_c4to2_sum_29_218, w_c4to2_carry_29_218, w_c4to2_cout_29_218;
math_compressor_4to2 u_c4to2_29_218 (
    .i_x1(w_c4to2_cout_28_114), .i_x2(w_c4to2_carry_28_115),
    .i_x3(w_c4to2_cout_28_115), .i_x4(w_c4to2_sum_29_116),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_218), .ow_carry(w_c4to2_carry_29_218), .ow_cout(w_c4to2_cout_29_218)
);
wire w_c4to2_sum_29_219, w_c4to2_carry_29_219, w_c4to2_cout_29_219;
math_compressor_4to2 u_c4to2_29_219 (
    .i_x1(w_c4to2_sum_29_117), .i_x2(w_c4to2_sum_29_118),
    .i_x3(w_c4to2_sum_29_119), .i_x4(w_c4to2_sum_29_120),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_219), .ow_carry(w_c4to2_carry_29_219), .ow_cout(w_c4to2_cout_29_219)
);
wire w_c4to2_sum_29_220, w_c4to2_carry_29_220, w_c4to2_cout_29_220;
math_compressor_4to2 u_c4to2_29_220 (
    .i_x1(w_c4to2_sum_29_121), .i_x2(w_c4to2_carry_28_213),
    .i_x3(w_c4to2_cout_28_213), .i_x4(w_c4to2_carry_28_214),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_220), .ow_carry(w_c4to2_carry_29_220), .ow_cout(w_c4to2_cout_29_220)
);
wire w_c4to2_sum_30_221, w_c4to2_carry_30_221, w_c4to2_cout_30_221;
math_compressor_4to2 u_c4to2_30_221 (
    .i_x1(w_c4to2_cout_29_118), .i_x2(w_c4to2_carry_29_119),
    .i_x3(w_c4to2_cout_29_119), .i_x4(w_c4to2_carry_29_120),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_221), .ow_carry(w_c4to2_carry_30_221), .ow_cout(w_c4to2_cout_30_221)
);
wire w_c4to2_sum_30_222, w_c4to2_carry_30_222, w_c4to2_cout_30_222;
math_compressor_4to2 u_c4to2_30_222 (
    .i_x1(w_c4to2_cout_29_120), .i_x2(w_c4to2_carry_29_121),
    .i_x3(w_c4to2_cout_29_121), .i_x4(w_c4to2_sum_30_122),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_222), .ow_carry(w_c4to2_carry_30_222), .ow_cout(w_c4to2_cout_30_222)
);
wire w_c4to2_sum_30_223, w_c4to2_carry_30_223, w_c4to2_cout_30_223;
math_compressor_4to2 u_c4to2_30_223 (
    .i_x1(w_c4to2_sum_30_123), .i_x2(w_c4to2_sum_30_124),
    .i_x3(w_c4to2_sum_30_125), .i_x4(w_c4to2_sum_30_126),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_223), .ow_carry(w_c4to2_carry_30_223), .ow_cout(w_c4to2_cout_30_223)
);
wire w_c4to2_sum_30_224, w_c4to2_carry_30_224, w_c4to2_cout_30_224;
math_compressor_4to2 u_c4to2_30_224 (
    .i_x1(w_c4to2_sum_30_127), .i_x2(w_c4to2_carry_29_217),
    .i_x3(w_c4to2_cout_29_217), .i_x4(w_c4to2_carry_29_218),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_224), .ow_carry(w_c4to2_carry_30_224), .ow_cout(w_c4to2_cout_30_224)
);
wire w_c4to2_sum_31_225, w_c4to2_carry_31_225, w_c4to2_cout_31_225;
math_compressor_4to2 u_c4to2_31_225 (
    .i_x1(w_c4to2_carry_30_124), .i_x2(w_c4to2_cout_30_124),
    .i_x3(w_c4to2_carry_30_125), .i_x4(w_c4to2_cout_30_125),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_225), .ow_carry(w_c4to2_carry_31_225), .ow_cout(w_c4to2_cout_31_225)
);
wire w_c4to2_sum_31_226, w_c4to2_carry_31_226, w_c4to2_cout_31_226;
math_compressor_4to2 u_c4to2_31_226 (
    .i_x1(w_c4to2_carry_30_126), .i_x2(w_c4to2_cout_30_126),
    .i_x3(w_c4to2_carry_30_127), .i_x4(w_c4to2_cout_30_127),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_226), .ow_carry(w_c4to2_carry_31_226), .ow_cout(w_c4to2_cout_31_226)
);
wire w_c4to2_sum_31_227, w_c4to2_carry_31_227, w_c4to2_cout_31_227;
math_compressor_4to2 u_c4to2_31_227 (
    .i_x1(w_c4to2_sum_31_128), .i_x2(w_c4to2_sum_31_129),
    .i_x3(w_c4to2_sum_31_130), .i_x4(w_c4to2_sum_31_131),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_227), .ow_carry(w_c4to2_carry_31_227), .ow_cout(w_c4to2_cout_31_227)
);
wire w_c4to2_sum_31_228, w_c4to2_carry_31_228, w_c4to2_cout_31_228;
math_compressor_4to2 u_c4to2_31_228 (
    .i_x1(w_c4to2_sum_31_132), .i_x2(w_c4to2_carry_30_221),
    .i_x3(w_c4to2_cout_30_221), .i_x4(w_c4to2_carry_30_222),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_228), .ow_carry(w_c4to2_carry_31_228), .ow_cout(w_c4to2_cout_31_228)
);
wire w_c4to2_sum_32_229, w_c4to2_carry_32_229, w_c4to2_cout_32_229;
math_compressor_4to2 u_c4to2_32_229 (
    .i_x1(w_c4to2_cout_31_128), .i_x2(w_c4to2_carry_31_129),
    .i_x3(w_c4to2_cout_31_129), .i_x4(w_c4to2_carry_31_130),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_229), .ow_carry(w_c4to2_carry_32_229), .ow_cout(w_c4to2_cout_32_229)
);
wire w_c4to2_sum_32_230, w_c4to2_carry_32_230, w_c4to2_cout_32_230;
math_compressor_4to2 u_c4to2_32_230 (
    .i_x1(w_c4to2_cout_31_130), .i_x2(w_c4to2_carry_31_131),
    .i_x3(w_c4to2_cout_31_131), .i_x4(w_c4to2_carry_31_132),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_230), .ow_carry(w_c4to2_carry_32_230), .ow_cout(w_c4to2_cout_32_230)
);
wire w_c4to2_sum_32_231, w_c4to2_carry_32_231, w_c4to2_cout_32_231;
math_compressor_4to2 u_c4to2_32_231 (
    .i_x1(w_c4to2_cout_31_132), .i_x2(w_c4to2_sum_32_133),
    .i_x3(w_c4to2_sum_32_134), .i_x4(w_c4to2_sum_32_135),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_231), .ow_carry(w_c4to2_carry_32_231), .ow_cout(w_c4to2_cout_32_231)
);
wire w_c4to2_sum_32_232, w_c4to2_carry_32_232, w_c4to2_cout_32_232;
math_compressor_4to2 u_c4to2_32_232 (
    .i_x1(w_c4to2_sum_32_136), .i_x2(w_c4to2_carry_31_225),
    .i_x3(w_c4to2_cout_31_225), .i_x4(w_c4to2_carry_31_226),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_232), .ow_carry(w_c4to2_carry_32_232), .ow_cout(w_c4to2_cout_32_232)
);
wire w_c4to2_sum_33_233, w_c4to2_carry_33_233, w_c4to2_cout_33_233;
math_compressor_4to2 u_c4to2_33_233 (
    .i_x1(w_pp_22_11), .i_x2(w_pp_23_10),
    .i_x3(w_c4to2_carry_32_133), .i_x4(w_c4to2_cout_32_133),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_233), .ow_carry(w_c4to2_carry_33_233), .ow_cout(w_c4to2_cout_33_233)
);
wire w_c4to2_sum_33_234, w_c4to2_carry_33_234, w_c4to2_cout_33_234;
math_compressor_4to2 u_c4to2_33_234 (
    .i_x1(w_c4to2_carry_32_134), .i_x2(w_c4to2_cout_32_134),
    .i_x3(w_c4to2_carry_32_135), .i_x4(w_c4to2_cout_32_135),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_234), .ow_carry(w_c4to2_carry_33_234), .ow_cout(w_c4to2_cout_33_234)
);
wire w_c4to2_sum_33_235, w_c4to2_carry_33_235, w_c4to2_cout_33_235;
math_compressor_4to2 u_c4to2_33_235 (
    .i_x1(w_c4to2_carry_32_136), .i_x2(w_c4to2_cout_32_136),
    .i_x3(w_c4to2_sum_33_137), .i_x4(w_c4to2_sum_33_138),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_235), .ow_carry(w_c4to2_carry_33_235), .ow_cout(w_c4to2_cout_33_235)
);
wire w_c4to2_sum_33_236, w_c4to2_carry_33_236, w_c4to2_cout_33_236;
math_compressor_4to2 u_c4to2_33_236 (
    .i_x1(w_c4to2_sum_33_139), .i_x2(w_c4to2_carry_32_229),
    .i_x3(w_c4to2_cout_32_229), .i_x4(w_c4to2_carry_32_230),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_236), .ow_carry(w_c4to2_carry_33_236), .ow_cout(w_c4to2_cout_33_236)
);
wire w_c4to2_sum_34_237, w_c4to2_carry_34_237, w_c4to2_cout_34_237;
math_compressor_4to2 u_c4to2_34_237 (
    .i_x1(w_pp_19_15), .i_x2(w_pp_20_14),
    .i_x3(w_pp_21_13), .i_x4(w_pp_22_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_237), .ow_carry(w_c4to2_carry_34_237), .ow_cout(w_c4to2_cout_34_237)
);
wire w_c4to2_sum_34_238, w_c4to2_carry_34_238, w_c4to2_cout_34_238;
math_compressor_4to2 u_c4to2_34_238 (
    .i_x1(w_pp_23_11), .i_x2(w_c4to2_carry_33_137),
    .i_x3(w_c4to2_cout_33_137), .i_x4(w_c4to2_carry_33_138),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_238), .ow_carry(w_c4to2_carry_34_238), .ow_cout(w_c4to2_cout_34_238)
);
wire w_c4to2_sum_34_239, w_c4to2_carry_34_239, w_c4to2_cout_34_239;
math_compressor_4to2 u_c4to2_34_239 (
    .i_x1(w_c4to2_cout_33_138), .i_x2(w_c4to2_carry_33_139),
    .i_x3(w_c4to2_cout_33_139), .i_x4(w_c4to2_sum_34_140),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_239), .ow_carry(w_c4to2_carry_34_239), .ow_cout(w_c4to2_cout_34_239)
);
wire w_c4to2_sum_34_240, w_c4to2_carry_34_240, w_c4to2_cout_34_240;
math_compressor_4to2 u_c4to2_34_240 (
    .i_x1(w_c4to2_sum_34_141), .i_x2(w_c4to2_carry_33_233),
    .i_x3(w_c4to2_cout_33_233), .i_x4(w_c4to2_carry_33_234),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_240), .ow_carry(w_c4to2_carry_34_240), .ow_cout(w_c4to2_cout_34_240)
);
wire w_c4to2_sum_35_241, w_c4to2_carry_35_241, w_c4to2_cout_35_241;
math_compressor_4to2 u_c4to2_35_241 (
    .i_x1(w_pp_16_19), .i_x2(w_pp_17_18),
    .i_x3(w_pp_18_17), .i_x4(w_pp_19_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_241), .ow_carry(w_c4to2_carry_35_241), .ow_cout(w_c4to2_cout_35_241)
);
wire w_c4to2_sum_35_242, w_c4to2_carry_35_242, w_c4to2_cout_35_242;
math_compressor_4to2 u_c4to2_35_242 (
    .i_x1(w_pp_20_15), .i_x2(w_pp_21_14),
    .i_x3(w_pp_22_13), .i_x4(w_pp_23_12),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_242), .ow_carry(w_c4to2_carry_35_242), .ow_cout(w_c4to2_cout_35_242)
);
wire w_c4to2_sum_35_243, w_c4to2_carry_35_243, w_c4to2_cout_35_243;
math_compressor_4to2 u_c4to2_35_243 (
    .i_x1(w_c4to2_carry_34_140), .i_x2(w_c4to2_cout_34_140),
    .i_x3(w_c4to2_carry_34_141), .i_x4(w_c4to2_cout_34_141),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_243), .ow_carry(w_c4to2_carry_35_243), .ow_cout(w_c4to2_cout_35_243)
);
wire w_c4to2_sum_35_244, w_c4to2_carry_35_244, w_c4to2_cout_35_244;
math_compressor_4to2 u_c4to2_35_244 (
    .i_x1(w_c4to2_sum_35_142), .i_x2(w_c4to2_carry_34_237),
    .i_x3(w_c4to2_cout_34_237), .i_x4(w_c4to2_carry_34_238),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_244), .ow_carry(w_c4to2_carry_35_244), .ow_cout(w_c4to2_cout_35_244)
);
wire w_c4to2_sum_36_245, w_c4to2_carry_36_245, w_c4to2_cout_36_245;
math_compressor_4to2 u_c4to2_36_245 (
    .i_x1(w_pp_13_23), .i_x2(w_pp_14_22),
    .i_x3(w_pp_15_21), .i_x4(w_pp_16_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_245), .ow_carry(w_c4to2_carry_36_245), .ow_cout(w_c4to2_cout_36_245)
);
wire w_c4to2_sum_36_246, w_c4to2_carry_36_246, w_c4to2_cout_36_246;
math_compressor_4to2 u_c4to2_36_246 (
    .i_x1(w_pp_17_19), .i_x2(w_pp_18_18),
    .i_x3(w_pp_19_17), .i_x4(w_pp_20_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_246), .ow_carry(w_c4to2_carry_36_246), .ow_cout(w_c4to2_cout_36_246)
);
wire w_c4to2_sum_36_247, w_c4to2_carry_36_247, w_c4to2_cout_36_247;
math_compressor_4to2 u_c4to2_36_247 (
    .i_x1(w_pp_21_15), .i_x2(w_pp_22_14),
    .i_x3(w_pp_23_13), .i_x4(w_c4to2_carry_35_142),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_247), .ow_carry(w_c4to2_carry_36_247), .ow_cout(w_c4to2_cout_36_247)
);
wire w_c4to2_sum_36_248, w_c4to2_carry_36_248, w_c4to2_cout_36_248;
math_compressor_4to2 u_c4to2_36_248 (
    .i_x1(w_c4to2_cout_35_142), .i_x2(w_c4to2_carry_35_241),
    .i_x3(w_c4to2_cout_35_241), .i_x4(w_c4to2_carry_35_242),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_248), .ow_carry(w_c4to2_carry_36_248), .ow_cout(w_c4to2_cout_36_248)
);
wire w_c4to2_sum_37_249, w_c4to2_carry_37_249, w_c4to2_cout_37_249;
math_compressor_4to2 u_c4to2_37_249 (
    .i_x1(w_pp_14_23), .i_x2(w_pp_15_22),
    .i_x3(w_pp_16_21), .i_x4(w_pp_17_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_249), .ow_carry(w_c4to2_carry_37_249), .ow_cout(w_c4to2_cout_37_249)
);
wire w_c4to2_sum_37_250, w_c4to2_carry_37_250, w_c4to2_cout_37_250;
math_compressor_4to2 u_c4to2_37_250 (
    .i_x1(w_pp_18_19), .i_x2(w_pp_19_18),
    .i_x3(w_pp_20_17), .i_x4(w_pp_21_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_250), .ow_carry(w_c4to2_carry_37_250), .ow_cout(w_c4to2_cout_37_250)
);
wire w_c4to2_sum_37_251, w_c4to2_carry_37_251, w_c4to2_cout_37_251;
math_compressor_4to2 u_c4to2_37_251 (
    .i_x1(w_pp_22_15), .i_x2(w_pp_23_14),
    .i_x3(w_c4to2_carry_36_245), .i_x4(w_c4to2_cout_36_245),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_251), .ow_carry(w_c4to2_carry_37_251), .ow_cout(w_c4to2_cout_37_251)
);
wire w_c4to2_sum_38_252, w_c4to2_carry_38_252, w_c4to2_cout_38_252;
math_compressor_4to2 u_c4to2_38_252 (
    .i_x1(w_pp_15_23), .i_x2(w_pp_16_22),
    .i_x3(w_pp_17_21), .i_x4(w_pp_18_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_252), .ow_carry(w_c4to2_carry_38_252), .ow_cout(w_c4to2_cout_38_252)
);
wire w_c4to2_sum_38_253, w_c4to2_carry_38_253, w_c4to2_cout_38_253;
math_compressor_4to2 u_c4to2_38_253 (
    .i_x1(w_pp_19_19), .i_x2(w_pp_20_18),
    .i_x3(w_pp_21_17), .i_x4(w_pp_22_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_253), .ow_carry(w_c4to2_carry_38_253), .ow_cout(w_c4to2_cout_38_253)
);
wire w_c4to2_sum_39_254, w_c4to2_carry_39_254, w_c4to2_cout_39_254;
math_compressor_4to2 u_c4to2_39_254 (
    .i_x1(w_pp_16_23), .i_x2(w_pp_17_22),
    .i_x3(w_pp_18_21), .i_x4(w_pp_19_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_254), .ow_carry(w_c4to2_carry_39_254), .ow_cout(w_c4to2_cout_39_254)
);

// Dadda Reduction Stage 4: height 9 -> 6

wire w_c4to2_sum_06_255, w_c4to2_carry_06_255, w_c4to2_cout_06_255;
math_compressor_4to2 u_c4to2_06_255 (
    .i_x1(w_pp_00_06), .i_x2(w_pp_01_05),
    .i_x3(w_pp_02_04), .i_x4(w_pp_03_03),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_06_255), .ow_carry(w_c4to2_carry_06_255), .ow_cout(w_c4to2_cout_06_255)
);
wire w_c4to2_sum_07_256, w_c4to2_carry_07_256, w_c4to2_cout_07_256;
math_compressor_4to2 u_c4to2_07_256 (
    .i_x1(w_pp_00_07), .i_x2(w_pp_01_06),
    .i_x3(w_pp_02_05), .i_x4(w_pp_03_04),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_07_256), .ow_carry(w_c4to2_carry_07_256), .ow_cout(w_c4to2_cout_07_256)
);
wire w_c4to2_sum_07_257, w_c4to2_carry_07_257, w_c4to2_cout_07_257;
math_compressor_4to2 u_c4to2_07_257 (
    .i_x1(w_pp_04_03), .i_x2(w_pp_05_02),
    .i_x3(w_pp_06_01), .i_x4(w_pp_07_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_07_257), .ow_carry(w_c4to2_carry_07_257), .ow_cout(w_c4to2_cout_07_257)
);
wire w_c4to2_sum_08_258, w_c4to2_carry_08_258, w_c4to2_cout_08_258;
math_compressor_4to2 u_c4to2_08_258 (
    .i_x1(w_pp_00_08), .i_x2(w_pp_01_07),
    .i_x3(w_pp_02_06), .i_x4(w_pp_03_05),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_258), .ow_carry(w_c4to2_carry_08_258), .ow_cout(w_c4to2_cout_08_258)
);
wire w_c4to2_sum_08_259, w_c4to2_carry_08_259, w_c4to2_cout_08_259;
math_compressor_4to2 u_c4to2_08_259 (
    .i_x1(w_pp_04_04), .i_x2(w_pp_05_03),
    .i_x3(w_pp_06_02), .i_x4(w_pp_07_01),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_259), .ow_carry(w_c4to2_carry_08_259), .ow_cout(w_c4to2_cout_08_259)
);
wire w_c4to2_sum_08_260, w_c4to2_carry_08_260, w_c4to2_cout_08_260;
math_compressor_4to2 u_c4to2_08_260 (
    .i_x1(w_pp_08_00), .i_x2(w_c4to2_carry_07_256),
    .i_x3(w_c4to2_cout_07_256), .i_x4(w_c4to2_carry_07_257),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_260), .ow_carry(w_c4to2_carry_08_260), .ow_cout(w_c4to2_cout_08_260)
);
wire w_c4to2_sum_09_261, w_c4to2_carry_09_261, w_c4to2_cout_09_261;
math_compressor_4to2 u_c4to2_09_261 (
    .i_x1(w_pp_04_05), .i_x2(w_pp_05_04),
    .i_x3(w_pp_06_03), .i_x4(w_pp_07_02),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_261), .ow_carry(w_c4to2_carry_09_261), .ow_cout(w_c4to2_cout_09_261)
);
wire w_c4to2_sum_09_262, w_c4to2_carry_09_262, w_c4to2_cout_09_262;
math_compressor_4to2 u_c4to2_09_262 (
    .i_x1(w_pp_08_01), .i_x2(w_pp_09_00),
    .i_x3(w_c4to2_sum_09_143), .i_x4(w_c4to2_carry_08_258),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_262), .ow_carry(w_c4to2_carry_09_262), .ow_cout(w_c4to2_cout_09_262)
);
wire w_c4to2_sum_09_263, w_c4to2_carry_09_263, w_c4to2_cout_09_263;
math_compressor_4to2 u_c4to2_09_263 (
    .i_x1(w_c4to2_cout_08_258), .i_x2(w_c4to2_carry_08_259),
    .i_x3(w_c4to2_cout_08_259), .i_x4(w_c4to2_carry_08_260),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_263), .ow_carry(w_c4to2_carry_09_263), .ow_cout(w_c4to2_cout_09_263)
);
wire w_c4to2_sum_10_264, w_c4to2_carry_10_264, w_c4to2_cout_10_264;
math_compressor_4to2 u_c4to2_10_264 (
    .i_x1(w_pp_08_02), .i_x2(w_pp_09_01),
    .i_x3(w_pp_10_00), .i_x4(w_c4to2_carry_09_143),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_264), .ow_carry(w_c4to2_carry_10_264), .ow_cout(w_c4to2_cout_10_264)
);
wire w_c4to2_sum_10_265, w_c4to2_carry_10_265, w_c4to2_cout_10_265;
math_compressor_4to2 u_c4to2_10_265 (
    .i_x1(w_c4to2_cout_09_143), .i_x2(w_c4to2_sum_10_144),
    .i_x3(w_c4to2_sum_10_145), .i_x4(w_c4to2_carry_09_261),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_265), .ow_carry(w_c4to2_carry_10_265), .ow_cout(w_c4to2_cout_10_265)
);
wire w_c4to2_sum_10_266, w_c4to2_carry_10_266, w_c4to2_cout_10_266;
math_compressor_4to2 u_c4to2_10_266 (
    .i_x1(w_c4to2_cout_09_261), .i_x2(w_c4to2_carry_09_262),
    .i_x3(w_c4to2_cout_09_262), .i_x4(w_c4to2_carry_09_263),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_266), .ow_carry(w_c4to2_carry_10_266), .ow_cout(w_c4to2_cout_10_266)
);
wire w_c4to2_sum_11_267, w_c4to2_carry_11_267, w_c4to2_cout_11_267;
math_compressor_4to2 u_c4to2_11_267 (
    .i_x1(w_c4to2_carry_10_144), .i_x2(w_c4to2_cout_10_144),
    .i_x3(w_c4to2_carry_10_145), .i_x4(w_c4to2_cout_10_145),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_267), .ow_carry(w_c4to2_carry_11_267), .ow_cout(w_c4to2_cout_11_267)
);
wire w_c4to2_sum_11_268, w_c4to2_carry_11_268, w_c4to2_cout_11_268;
math_compressor_4to2 u_c4to2_11_268 (
    .i_x1(w_c4to2_sum_11_146), .i_x2(w_c4to2_sum_11_147),
    .i_x3(w_c4to2_sum_11_148), .i_x4(w_c4to2_carry_10_264),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_268), .ow_carry(w_c4to2_carry_11_268), .ow_cout(w_c4to2_cout_11_268)
);
wire w_c4to2_sum_11_269, w_c4to2_carry_11_269, w_c4to2_cout_11_269;
math_compressor_4to2 u_c4to2_11_269 (
    .i_x1(w_c4to2_cout_10_264), .i_x2(w_c4to2_carry_10_265),
    .i_x3(w_c4to2_cout_10_265), .i_x4(w_c4to2_carry_10_266),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_269), .ow_carry(w_c4to2_carry_11_269), .ow_cout(w_c4to2_cout_11_269)
);
wire w_c4to2_sum_12_270, w_c4to2_carry_12_270, w_c4to2_cout_12_270;
math_compressor_4to2 u_c4to2_12_270 (
    .i_x1(w_c4to2_cout_11_147), .i_x2(w_c4to2_carry_11_148),
    .i_x3(w_c4to2_cout_11_148), .i_x4(w_c4to2_sum_12_149),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_270), .ow_carry(w_c4to2_carry_12_270), .ow_cout(w_c4to2_cout_12_270)
);
wire w_c4to2_sum_12_271, w_c4to2_carry_12_271, w_c4to2_cout_12_271;
math_compressor_4to2 u_c4to2_12_271 (
    .i_x1(w_c4to2_sum_12_150), .i_x2(w_c4to2_sum_12_151),
    .i_x3(w_c4to2_sum_12_152), .i_x4(w_c4to2_carry_11_267),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_271), .ow_carry(w_c4to2_carry_12_271), .ow_cout(w_c4to2_cout_12_271)
);
wire w_c4to2_sum_12_272, w_c4to2_carry_12_272, w_c4to2_cout_12_272;
math_compressor_4to2 u_c4to2_12_272 (
    .i_x1(w_c4to2_cout_11_267), .i_x2(w_c4to2_carry_11_268),
    .i_x3(w_c4to2_cout_11_268), .i_x4(w_c4to2_carry_11_269),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_272), .ow_carry(w_c4to2_carry_12_272), .ow_cout(w_c4to2_cout_12_272)
);
wire w_c4to2_sum_13_273, w_c4to2_carry_13_273, w_c4to2_cout_13_273;
math_compressor_4to2 u_c4to2_13_273 (
    .i_x1(w_c4to2_cout_12_151), .i_x2(w_c4to2_carry_12_152),
    .i_x3(w_c4to2_cout_12_152), .i_x4(w_c4to2_sum_13_153),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_273), .ow_carry(w_c4to2_carry_13_273), .ow_cout(w_c4to2_cout_13_273)
);
wire w_c4to2_sum_13_274, w_c4to2_carry_13_274, w_c4to2_cout_13_274;
math_compressor_4to2 u_c4to2_13_274 (
    .i_x1(w_c4to2_sum_13_154), .i_x2(w_c4to2_sum_13_155),
    .i_x3(w_c4to2_sum_13_156), .i_x4(w_c4to2_carry_12_270),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_274), .ow_carry(w_c4to2_carry_13_274), .ow_cout(w_c4to2_cout_13_274)
);
wire w_c4to2_sum_13_275, w_c4to2_carry_13_275, w_c4to2_cout_13_275;
math_compressor_4to2 u_c4to2_13_275 (
    .i_x1(w_c4to2_cout_12_270), .i_x2(w_c4to2_carry_12_271),
    .i_x3(w_c4to2_cout_12_271), .i_x4(w_c4to2_carry_12_272),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_275), .ow_carry(w_c4to2_carry_13_275), .ow_cout(w_c4to2_cout_13_275)
);
wire w_c4to2_sum_14_276, w_c4to2_carry_14_276, w_c4to2_cout_14_276;
math_compressor_4to2 u_c4to2_14_276 (
    .i_x1(w_c4to2_cout_13_155), .i_x2(w_c4to2_carry_13_156),
    .i_x3(w_c4to2_cout_13_156), .i_x4(w_c4to2_sum_14_157),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_276), .ow_carry(w_c4to2_carry_14_276), .ow_cout(w_c4to2_cout_14_276)
);
wire w_c4to2_sum_14_277, w_c4to2_carry_14_277, w_c4to2_cout_14_277;
math_compressor_4to2 u_c4to2_14_277 (
    .i_x1(w_c4to2_sum_14_158), .i_x2(w_c4to2_sum_14_159),
    .i_x3(w_c4to2_sum_14_160), .i_x4(w_c4to2_carry_13_273),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_277), .ow_carry(w_c4to2_carry_14_277), .ow_cout(w_c4to2_cout_14_277)
);
wire w_c4to2_sum_14_278, w_c4to2_carry_14_278, w_c4to2_cout_14_278;
math_compressor_4to2 u_c4to2_14_278 (
    .i_x1(w_c4to2_cout_13_273), .i_x2(w_c4to2_carry_13_274),
    .i_x3(w_c4to2_cout_13_274), .i_x4(w_c4to2_carry_13_275),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_278), .ow_carry(w_c4to2_carry_14_278), .ow_cout(w_c4to2_cout_14_278)
);
wire w_c4to2_sum_15_279, w_c4to2_carry_15_279, w_c4to2_cout_15_279;
math_compressor_4to2 u_c4to2_15_279 (
    .i_x1(w_c4to2_cout_14_159), .i_x2(w_c4to2_carry_14_160),
    .i_x3(w_c4to2_cout_14_160), .i_x4(w_c4to2_sum_15_161),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_279), .ow_carry(w_c4to2_carry_15_279), .ow_cout(w_c4to2_cout_15_279)
);
wire w_c4to2_sum_15_280, w_c4to2_carry_15_280, w_c4to2_cout_15_280;
math_compressor_4to2 u_c4to2_15_280 (
    .i_x1(w_c4to2_sum_15_162), .i_x2(w_c4to2_sum_15_163),
    .i_x3(w_c4to2_sum_15_164), .i_x4(w_c4to2_carry_14_276),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_280), .ow_carry(w_c4to2_carry_15_280), .ow_cout(w_c4to2_cout_15_280)
);
wire w_c4to2_sum_15_281, w_c4to2_carry_15_281, w_c4to2_cout_15_281;
math_compressor_4to2 u_c4to2_15_281 (
    .i_x1(w_c4to2_cout_14_276), .i_x2(w_c4to2_carry_14_277),
    .i_x3(w_c4to2_cout_14_277), .i_x4(w_c4to2_carry_14_278),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_281), .ow_carry(w_c4to2_carry_15_281), .ow_cout(w_c4to2_cout_15_281)
);
wire w_c4to2_sum_16_282, w_c4to2_carry_16_282, w_c4to2_cout_16_282;
math_compressor_4to2 u_c4to2_16_282 (
    .i_x1(w_c4to2_cout_15_163), .i_x2(w_c4to2_carry_15_164),
    .i_x3(w_c4to2_cout_15_164), .i_x4(w_c4to2_sum_16_165),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_282), .ow_carry(w_c4to2_carry_16_282), .ow_cout(w_c4to2_cout_16_282)
);
wire w_c4to2_sum_16_283, w_c4to2_carry_16_283, w_c4to2_cout_16_283;
math_compressor_4to2 u_c4to2_16_283 (
    .i_x1(w_c4to2_sum_16_166), .i_x2(w_c4to2_sum_16_167),
    .i_x3(w_c4to2_sum_16_168), .i_x4(w_c4to2_carry_15_279),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_283), .ow_carry(w_c4to2_carry_16_283), .ow_cout(w_c4to2_cout_16_283)
);
wire w_c4to2_sum_16_284, w_c4to2_carry_16_284, w_c4to2_cout_16_284;
math_compressor_4to2 u_c4to2_16_284 (
    .i_x1(w_c4to2_cout_15_279), .i_x2(w_c4to2_carry_15_280),
    .i_x3(w_c4to2_cout_15_280), .i_x4(w_c4to2_carry_15_281),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_284), .ow_carry(w_c4to2_carry_16_284), .ow_cout(w_c4to2_cout_16_284)
);
wire w_c4to2_sum_17_285, w_c4to2_carry_17_285, w_c4to2_cout_17_285;
math_compressor_4to2 u_c4to2_17_285 (
    .i_x1(w_c4to2_cout_16_167), .i_x2(w_c4to2_carry_16_168),
    .i_x3(w_c4to2_cout_16_168), .i_x4(w_c4to2_sum_17_169),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_285), .ow_carry(w_c4to2_carry_17_285), .ow_cout(w_c4to2_cout_17_285)
);
wire w_c4to2_sum_17_286, w_c4to2_carry_17_286, w_c4to2_cout_17_286;
math_compressor_4to2 u_c4to2_17_286 (
    .i_x1(w_c4to2_sum_17_170), .i_x2(w_c4to2_sum_17_171),
    .i_x3(w_c4to2_sum_17_172), .i_x4(w_c4to2_carry_16_282),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_286), .ow_carry(w_c4to2_carry_17_286), .ow_cout(w_c4to2_cout_17_286)
);
wire w_c4to2_sum_17_287, w_c4to2_carry_17_287, w_c4to2_cout_17_287;
math_compressor_4to2 u_c4to2_17_287 (
    .i_x1(w_c4to2_cout_16_282), .i_x2(w_c4to2_carry_16_283),
    .i_x3(w_c4to2_cout_16_283), .i_x4(w_c4to2_carry_16_284),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_287), .ow_carry(w_c4to2_carry_17_287), .ow_cout(w_c4to2_cout_17_287)
);
wire w_c4to2_sum_18_288, w_c4to2_carry_18_288, w_c4to2_cout_18_288;
math_compressor_4to2 u_c4to2_18_288 (
    .i_x1(w_c4to2_cout_17_171), .i_x2(w_c4to2_carry_17_172),
    .i_x3(w_c4to2_cout_17_172), .i_x4(w_c4to2_sum_18_173),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_288), .ow_carry(w_c4to2_carry_18_288), .ow_cout(w_c4to2_cout_18_288)
);
wire w_c4to2_sum_18_289, w_c4to2_carry_18_289, w_c4to2_cout_18_289;
math_compressor_4to2 u_c4to2_18_289 (
    .i_x1(w_c4to2_sum_18_174), .i_x2(w_c4to2_sum_18_175),
    .i_x3(w_c4to2_sum_18_176), .i_x4(w_c4to2_carry_17_285),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_289), .ow_carry(w_c4to2_carry_18_289), .ow_cout(w_c4to2_cout_18_289)
);
wire w_c4to2_sum_18_290, w_c4to2_carry_18_290, w_c4to2_cout_18_290;
math_compressor_4to2 u_c4to2_18_290 (
    .i_x1(w_c4to2_cout_17_285), .i_x2(w_c4to2_carry_17_286),
    .i_x3(w_c4to2_cout_17_286), .i_x4(w_c4to2_carry_17_287),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_290), .ow_carry(w_c4to2_carry_18_290), .ow_cout(w_c4to2_cout_18_290)
);
wire w_c4to2_sum_19_291, w_c4to2_carry_19_291, w_c4to2_cout_19_291;
math_compressor_4to2 u_c4to2_19_291 (
    .i_x1(w_c4to2_cout_18_175), .i_x2(w_c4to2_carry_18_176),
    .i_x3(w_c4to2_cout_18_176), .i_x4(w_c4to2_sum_19_177),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_291), .ow_carry(w_c4to2_carry_19_291), .ow_cout(w_c4to2_cout_19_291)
);
wire w_c4to2_sum_19_292, w_c4to2_carry_19_292, w_c4to2_cout_19_292;
math_compressor_4to2 u_c4to2_19_292 (
    .i_x1(w_c4to2_sum_19_178), .i_x2(w_c4to2_sum_19_179),
    .i_x3(w_c4to2_sum_19_180), .i_x4(w_c4to2_carry_18_288),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_292), .ow_carry(w_c4to2_carry_19_292), .ow_cout(w_c4to2_cout_19_292)
);
wire w_c4to2_sum_19_293, w_c4to2_carry_19_293, w_c4to2_cout_19_293;
math_compressor_4to2 u_c4to2_19_293 (
    .i_x1(w_c4to2_cout_18_288), .i_x2(w_c4to2_carry_18_289),
    .i_x3(w_c4to2_cout_18_289), .i_x4(w_c4to2_carry_18_290),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_293), .ow_carry(w_c4to2_carry_19_293), .ow_cout(w_c4to2_cout_19_293)
);
wire w_c4to2_sum_20_294, w_c4to2_carry_20_294, w_c4to2_cout_20_294;
math_compressor_4to2 u_c4to2_20_294 (
    .i_x1(w_c4to2_cout_19_179), .i_x2(w_c4to2_carry_19_180),
    .i_x3(w_c4to2_cout_19_180), .i_x4(w_c4to2_sum_20_181),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_294), .ow_carry(w_c4to2_carry_20_294), .ow_cout(w_c4to2_cout_20_294)
);
wire w_c4to2_sum_20_295, w_c4to2_carry_20_295, w_c4to2_cout_20_295;
math_compressor_4to2 u_c4to2_20_295 (
    .i_x1(w_c4to2_sum_20_182), .i_x2(w_c4to2_sum_20_183),
    .i_x3(w_c4to2_sum_20_184), .i_x4(w_c4to2_carry_19_291),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_295), .ow_carry(w_c4to2_carry_20_295), .ow_cout(w_c4to2_cout_20_295)
);
wire w_c4to2_sum_20_296, w_c4to2_carry_20_296, w_c4to2_cout_20_296;
math_compressor_4to2 u_c4to2_20_296 (
    .i_x1(w_c4to2_cout_19_291), .i_x2(w_c4to2_carry_19_292),
    .i_x3(w_c4to2_cout_19_292), .i_x4(w_c4to2_carry_19_293),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_296), .ow_carry(w_c4to2_carry_20_296), .ow_cout(w_c4to2_cout_20_296)
);
wire w_c4to2_sum_21_297, w_c4to2_carry_21_297, w_c4to2_cout_21_297;
math_compressor_4to2 u_c4to2_21_297 (
    .i_x1(w_c4to2_cout_20_183), .i_x2(w_c4to2_carry_20_184),
    .i_x3(w_c4to2_cout_20_184), .i_x4(w_c4to2_sum_21_185),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_297), .ow_carry(w_c4to2_carry_21_297), .ow_cout(w_c4to2_cout_21_297)
);
wire w_c4to2_sum_21_298, w_c4to2_carry_21_298, w_c4to2_cout_21_298;
math_compressor_4to2 u_c4to2_21_298 (
    .i_x1(w_c4to2_sum_21_186), .i_x2(w_c4to2_sum_21_187),
    .i_x3(w_c4to2_sum_21_188), .i_x4(w_c4to2_carry_20_294),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_298), .ow_carry(w_c4to2_carry_21_298), .ow_cout(w_c4to2_cout_21_298)
);
wire w_c4to2_sum_21_299, w_c4to2_carry_21_299, w_c4to2_cout_21_299;
math_compressor_4to2 u_c4to2_21_299 (
    .i_x1(w_c4to2_cout_20_294), .i_x2(w_c4to2_carry_20_295),
    .i_x3(w_c4to2_cout_20_295), .i_x4(w_c4to2_carry_20_296),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_299), .ow_carry(w_c4to2_carry_21_299), .ow_cout(w_c4to2_cout_21_299)
);
wire w_c4to2_sum_22_300, w_c4to2_carry_22_300, w_c4to2_cout_22_300;
math_compressor_4to2 u_c4to2_22_300 (
    .i_x1(w_c4to2_cout_21_187), .i_x2(w_c4to2_carry_21_188),
    .i_x3(w_c4to2_cout_21_188), .i_x4(w_c4to2_sum_22_189),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_300), .ow_carry(w_c4to2_carry_22_300), .ow_cout(w_c4to2_cout_22_300)
);
wire w_c4to2_sum_22_301, w_c4to2_carry_22_301, w_c4to2_cout_22_301;
math_compressor_4to2 u_c4to2_22_301 (
    .i_x1(w_c4to2_sum_22_190), .i_x2(w_c4to2_sum_22_191),
    .i_x3(w_c4to2_sum_22_192), .i_x4(w_c4to2_carry_21_297),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_301), .ow_carry(w_c4to2_carry_22_301), .ow_cout(w_c4to2_cout_22_301)
);
wire w_c4to2_sum_22_302, w_c4to2_carry_22_302, w_c4to2_cout_22_302;
math_compressor_4to2 u_c4to2_22_302 (
    .i_x1(w_c4to2_cout_21_297), .i_x2(w_c4to2_carry_21_298),
    .i_x3(w_c4to2_cout_21_298), .i_x4(w_c4to2_carry_21_299),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_302), .ow_carry(w_c4to2_carry_22_302), .ow_cout(w_c4to2_cout_22_302)
);
wire w_c4to2_sum_23_303, w_c4to2_carry_23_303, w_c4to2_cout_23_303;
math_compressor_4to2 u_c4to2_23_303 (
    .i_x1(w_c4to2_cout_22_191), .i_x2(w_c4to2_carry_22_192),
    .i_x3(w_c4to2_cout_22_192), .i_x4(w_c4to2_sum_23_193),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_303), .ow_carry(w_c4to2_carry_23_303), .ow_cout(w_c4to2_cout_23_303)
);
wire w_c4to2_sum_23_304, w_c4to2_carry_23_304, w_c4to2_cout_23_304;
math_compressor_4to2 u_c4to2_23_304 (
    .i_x1(w_c4to2_sum_23_194), .i_x2(w_c4to2_sum_23_195),
    .i_x3(w_c4to2_sum_23_196), .i_x4(w_c4to2_carry_22_300),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_304), .ow_carry(w_c4to2_carry_23_304), .ow_cout(w_c4to2_cout_23_304)
);
wire w_c4to2_sum_23_305, w_c4to2_carry_23_305, w_c4to2_cout_23_305;
math_compressor_4to2 u_c4to2_23_305 (
    .i_x1(w_c4to2_cout_22_300), .i_x2(w_c4to2_carry_22_301),
    .i_x3(w_c4to2_cout_22_301), .i_x4(w_c4to2_carry_22_302),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_305), .ow_carry(w_c4to2_carry_23_305), .ow_cout(w_c4to2_cout_23_305)
);
wire w_c4to2_sum_24_306, w_c4to2_carry_24_306, w_c4to2_cout_24_306;
math_compressor_4to2 u_c4to2_24_306 (
    .i_x1(w_c4to2_carry_23_195), .i_x2(w_c4to2_cout_23_195),
    .i_x3(w_c4to2_carry_23_196), .i_x4(w_c4to2_cout_23_196),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_306), .ow_carry(w_c4to2_carry_24_306), .ow_cout(w_c4to2_cout_24_306)
);
wire w_c4to2_sum_24_307, w_c4to2_carry_24_307, w_c4to2_cout_24_307;
math_compressor_4to2 u_c4to2_24_307 (
    .i_x1(w_c4to2_sum_24_197), .i_x2(w_c4to2_sum_24_198),
    .i_x3(w_c4to2_sum_24_199), .i_x4(w_c4to2_sum_24_200),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_307), .ow_carry(w_c4to2_carry_24_307), .ow_cout(w_c4to2_cout_24_307)
);
wire w_c4to2_sum_24_308, w_c4to2_carry_24_308, w_c4to2_cout_24_308;
math_compressor_4to2 u_c4to2_24_308 (
    .i_x1(w_c4to2_carry_23_303), .i_x2(w_c4to2_cout_23_303),
    .i_x3(w_c4to2_carry_23_304), .i_x4(w_c4to2_cout_23_304),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_308), .ow_carry(w_c4to2_carry_24_308), .ow_cout(w_c4to2_cout_24_308)
);
wire w_c4to2_sum_25_309, w_c4to2_carry_25_309, w_c4to2_cout_25_309;
math_compressor_4to2 u_c4to2_25_309 (
    .i_x1(w_c4to2_cout_24_199), .i_x2(w_c4to2_carry_24_200),
    .i_x3(w_c4to2_cout_24_200), .i_x4(w_c4to2_sum_25_201),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_309), .ow_carry(w_c4to2_carry_25_309), .ow_cout(w_c4to2_cout_25_309)
);
wire w_c4to2_sum_25_310, w_c4to2_carry_25_310, w_c4to2_cout_25_310;
math_compressor_4to2 u_c4to2_25_310 (
    .i_x1(w_c4to2_sum_25_202), .i_x2(w_c4to2_sum_25_203),
    .i_x3(w_c4to2_sum_25_204), .i_x4(w_c4to2_carry_24_306),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_310), .ow_carry(w_c4to2_carry_25_310), .ow_cout(w_c4to2_cout_25_310)
);
wire w_c4to2_sum_25_311, w_c4to2_carry_25_311, w_c4to2_cout_25_311;
math_compressor_4to2 u_c4to2_25_311 (
    .i_x1(w_c4to2_cout_24_306), .i_x2(w_c4to2_carry_24_307),
    .i_x3(w_c4to2_cout_24_307), .i_x4(w_c4to2_carry_24_308),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_311), .ow_carry(w_c4to2_carry_25_311), .ow_cout(w_c4to2_cout_25_311)
);
wire w_c4to2_sum_26_312, w_c4to2_carry_26_312, w_c4to2_cout_26_312;
math_compressor_4to2 u_c4to2_26_312 (
    .i_x1(w_c4to2_cout_25_202), .i_x2(w_c4to2_carry_25_203),
    .i_x3(w_c4to2_cout_25_203), .i_x4(w_c4to2_carry_25_204),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_312), .ow_carry(w_c4to2_carry_26_312), .ow_cout(w_c4to2_cout_26_312)
);
wire w_c4to2_sum_26_313, w_c4to2_carry_26_313, w_c4to2_cout_26_313;
math_compressor_4to2 u_c4to2_26_313 (
    .i_x1(w_c4to2_cout_25_204), .i_x2(w_c4to2_sum_26_205),
    .i_x3(w_c4to2_sum_26_206), .i_x4(w_c4to2_sum_26_207),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_313), .ow_carry(w_c4to2_carry_26_313), .ow_cout(w_c4to2_cout_26_313)
);
wire w_c4to2_sum_26_314, w_c4to2_carry_26_314, w_c4to2_cout_26_314;
math_compressor_4to2 u_c4to2_26_314 (
    .i_x1(w_c4to2_sum_26_208), .i_x2(w_c4to2_carry_25_309),
    .i_x3(w_c4to2_cout_25_309), .i_x4(w_c4to2_carry_25_310),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_314), .ow_carry(w_c4to2_carry_26_314), .ow_cout(w_c4to2_cout_26_314)
);
wire w_c4to2_sum_27_315, w_c4to2_carry_27_315, w_c4to2_cout_27_315;
math_compressor_4to2 u_c4to2_27_315 (
    .i_x1(w_c4to2_cout_26_206), .i_x2(w_c4to2_carry_26_207),
    .i_x3(w_c4to2_cout_26_207), .i_x4(w_c4to2_carry_26_208),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_315), .ow_carry(w_c4to2_carry_27_315), .ow_cout(w_c4to2_cout_27_315)
);
wire w_c4to2_sum_27_316, w_c4to2_carry_27_316, w_c4to2_cout_27_316;
math_compressor_4to2 u_c4to2_27_316 (
    .i_x1(w_c4to2_cout_26_208), .i_x2(w_c4to2_sum_27_209),
    .i_x3(w_c4to2_sum_27_210), .i_x4(w_c4to2_sum_27_211),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_316), .ow_carry(w_c4to2_carry_27_316), .ow_cout(w_c4to2_cout_27_316)
);
wire w_c4to2_sum_27_317, w_c4to2_carry_27_317, w_c4to2_cout_27_317;
math_compressor_4to2 u_c4to2_27_317 (
    .i_x1(w_c4to2_sum_27_212), .i_x2(w_c4to2_carry_26_312),
    .i_x3(w_c4to2_cout_26_312), .i_x4(w_c4to2_carry_26_313),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_317), .ow_carry(w_c4to2_carry_27_317), .ow_cout(w_c4to2_cout_27_317)
);
wire w_c4to2_sum_28_318, w_c4to2_carry_28_318, w_c4to2_cout_28_318;
math_compressor_4to2 u_c4to2_28_318 (
    .i_x1(w_c4to2_cout_27_210), .i_x2(w_c4to2_carry_27_211),
    .i_x3(w_c4to2_cout_27_211), .i_x4(w_c4to2_carry_27_212),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_318), .ow_carry(w_c4to2_carry_28_318), .ow_cout(w_c4to2_cout_28_318)
);
wire w_c4to2_sum_28_319, w_c4to2_carry_28_319, w_c4to2_cout_28_319;
math_compressor_4to2 u_c4to2_28_319 (
    .i_x1(w_c4to2_cout_27_212), .i_x2(w_c4to2_sum_28_213),
    .i_x3(w_c4to2_sum_28_214), .i_x4(w_c4to2_sum_28_215),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_319), .ow_carry(w_c4to2_carry_28_319), .ow_cout(w_c4to2_cout_28_319)
);
wire w_c4to2_sum_28_320, w_c4to2_carry_28_320, w_c4to2_cout_28_320;
math_compressor_4to2 u_c4to2_28_320 (
    .i_x1(w_c4to2_sum_28_216), .i_x2(w_c4to2_carry_27_315),
    .i_x3(w_c4to2_cout_27_315), .i_x4(w_c4to2_carry_27_316),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_320), .ow_carry(w_c4to2_carry_28_320), .ow_cout(w_c4to2_cout_28_320)
);
wire w_c4to2_sum_29_321, w_c4to2_carry_29_321, w_c4to2_cout_29_321;
math_compressor_4to2 u_c4to2_29_321 (
    .i_x1(w_c4to2_cout_28_214), .i_x2(w_c4to2_carry_28_215),
    .i_x3(w_c4to2_cout_28_215), .i_x4(w_c4to2_carry_28_216),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_321), .ow_carry(w_c4to2_carry_29_321), .ow_cout(w_c4to2_cout_29_321)
);
wire w_c4to2_sum_29_322, w_c4to2_carry_29_322, w_c4to2_cout_29_322;
math_compressor_4to2 u_c4to2_29_322 (
    .i_x1(w_c4to2_cout_28_216), .i_x2(w_c4to2_sum_29_217),
    .i_x3(w_c4to2_sum_29_218), .i_x4(w_c4to2_sum_29_219),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_322), .ow_carry(w_c4to2_carry_29_322), .ow_cout(w_c4to2_cout_29_322)
);
wire w_c4to2_sum_29_323, w_c4to2_carry_29_323, w_c4to2_cout_29_323;
math_compressor_4to2 u_c4to2_29_323 (
    .i_x1(w_c4to2_sum_29_220), .i_x2(w_c4to2_carry_28_318),
    .i_x3(w_c4to2_cout_28_318), .i_x4(w_c4to2_carry_28_319),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_323), .ow_carry(w_c4to2_carry_29_323), .ow_cout(w_c4to2_cout_29_323)
);
wire w_c4to2_sum_30_324, w_c4to2_carry_30_324, w_c4to2_cout_30_324;
math_compressor_4to2 u_c4to2_30_324 (
    .i_x1(w_c4to2_cout_29_218), .i_x2(w_c4to2_carry_29_219),
    .i_x3(w_c4to2_cout_29_219), .i_x4(w_c4to2_carry_29_220),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_324), .ow_carry(w_c4to2_carry_30_324), .ow_cout(w_c4to2_cout_30_324)
);
wire w_c4to2_sum_30_325, w_c4to2_carry_30_325, w_c4to2_cout_30_325;
math_compressor_4to2 u_c4to2_30_325 (
    .i_x1(w_c4to2_cout_29_220), .i_x2(w_c4to2_sum_30_221),
    .i_x3(w_c4to2_sum_30_222), .i_x4(w_c4to2_sum_30_223),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_325), .ow_carry(w_c4to2_carry_30_325), .ow_cout(w_c4to2_cout_30_325)
);
wire w_c4to2_sum_30_326, w_c4to2_carry_30_326, w_c4to2_cout_30_326;
math_compressor_4to2 u_c4to2_30_326 (
    .i_x1(w_c4to2_sum_30_224), .i_x2(w_c4to2_carry_29_321),
    .i_x3(w_c4to2_cout_29_321), .i_x4(w_c4to2_carry_29_322),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_326), .ow_carry(w_c4to2_carry_30_326), .ow_cout(w_c4to2_cout_30_326)
);
wire w_c4to2_sum_31_327, w_c4to2_carry_31_327, w_c4to2_cout_31_327;
math_compressor_4to2 u_c4to2_31_327 (
    .i_x1(w_c4to2_cout_30_222), .i_x2(w_c4to2_carry_30_223),
    .i_x3(w_c4to2_cout_30_223), .i_x4(w_c4to2_carry_30_224),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_327), .ow_carry(w_c4to2_carry_31_327), .ow_cout(w_c4to2_cout_31_327)
);
wire w_c4to2_sum_31_328, w_c4to2_carry_31_328, w_c4to2_cout_31_328;
math_compressor_4to2 u_c4to2_31_328 (
    .i_x1(w_c4to2_cout_30_224), .i_x2(w_c4to2_sum_31_225),
    .i_x3(w_c4to2_sum_31_226), .i_x4(w_c4to2_sum_31_227),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_328), .ow_carry(w_c4to2_carry_31_328), .ow_cout(w_c4to2_cout_31_328)
);
wire w_c4to2_sum_31_329, w_c4to2_carry_31_329, w_c4to2_cout_31_329;
math_compressor_4to2 u_c4to2_31_329 (
    .i_x1(w_c4to2_sum_31_228), .i_x2(w_c4to2_carry_30_324),
    .i_x3(w_c4to2_cout_30_324), .i_x4(w_c4to2_carry_30_325),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_329), .ow_carry(w_c4to2_carry_31_329), .ow_cout(w_c4to2_cout_31_329)
);
wire w_c4to2_sum_32_330, w_c4to2_carry_32_330, w_c4to2_cout_32_330;
math_compressor_4to2 u_c4to2_32_330 (
    .i_x1(w_c4to2_cout_31_226), .i_x2(w_c4to2_carry_31_227),
    .i_x3(w_c4to2_cout_31_227), .i_x4(w_c4to2_carry_31_228),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_330), .ow_carry(w_c4to2_carry_32_330), .ow_cout(w_c4to2_cout_32_330)
);
wire w_c4to2_sum_32_331, w_c4to2_carry_32_331, w_c4to2_cout_32_331;
math_compressor_4to2 u_c4to2_32_331 (
    .i_x1(w_c4to2_cout_31_228), .i_x2(w_c4to2_sum_32_229),
    .i_x3(w_c4to2_sum_32_230), .i_x4(w_c4to2_sum_32_231),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_331), .ow_carry(w_c4to2_carry_32_331), .ow_cout(w_c4to2_cout_32_331)
);
wire w_c4to2_sum_32_332, w_c4to2_carry_32_332, w_c4to2_cout_32_332;
math_compressor_4to2 u_c4to2_32_332 (
    .i_x1(w_c4to2_sum_32_232), .i_x2(w_c4to2_carry_31_327),
    .i_x3(w_c4to2_cout_31_327), .i_x4(w_c4to2_carry_31_328),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_332), .ow_carry(w_c4to2_carry_32_332), .ow_cout(w_c4to2_cout_32_332)
);
wire w_c4to2_sum_33_333, w_c4to2_carry_33_333, w_c4to2_cout_33_333;
math_compressor_4to2 u_c4to2_33_333 (
    .i_x1(w_c4to2_cout_32_230), .i_x2(w_c4to2_carry_32_231),
    .i_x3(w_c4to2_cout_32_231), .i_x4(w_c4to2_carry_32_232),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_333), .ow_carry(w_c4to2_carry_33_333), .ow_cout(w_c4to2_cout_33_333)
);
wire w_c4to2_sum_33_334, w_c4to2_carry_33_334, w_c4to2_cout_33_334;
math_compressor_4to2 u_c4to2_33_334 (
    .i_x1(w_c4to2_cout_32_232), .i_x2(w_c4to2_sum_33_233),
    .i_x3(w_c4to2_sum_33_234), .i_x4(w_c4to2_sum_33_235),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_334), .ow_carry(w_c4to2_carry_33_334), .ow_cout(w_c4to2_cout_33_334)
);
wire w_c4to2_sum_33_335, w_c4to2_carry_33_335, w_c4to2_cout_33_335;
math_compressor_4to2 u_c4to2_33_335 (
    .i_x1(w_c4to2_sum_33_236), .i_x2(w_c4to2_carry_32_330),
    .i_x3(w_c4to2_cout_32_330), .i_x4(w_c4to2_carry_32_331),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_335), .ow_carry(w_c4to2_carry_33_335), .ow_cout(w_c4to2_cout_33_335)
);
wire w_c4to2_sum_34_336, w_c4to2_carry_34_336, w_c4to2_cout_34_336;
math_compressor_4to2 u_c4to2_34_336 (
    .i_x1(w_c4to2_cout_33_234), .i_x2(w_c4to2_carry_33_235),
    .i_x3(w_c4to2_cout_33_235), .i_x4(w_c4to2_carry_33_236),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_336), .ow_carry(w_c4to2_carry_34_336), .ow_cout(w_c4to2_cout_34_336)
);
wire w_c4to2_sum_34_337, w_c4to2_carry_34_337, w_c4to2_cout_34_337;
math_compressor_4to2 u_c4to2_34_337 (
    .i_x1(w_c4to2_cout_33_236), .i_x2(w_c4to2_sum_34_237),
    .i_x3(w_c4to2_sum_34_238), .i_x4(w_c4to2_sum_34_239),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_337), .ow_carry(w_c4to2_carry_34_337), .ow_cout(w_c4to2_cout_34_337)
);
wire w_c4to2_sum_34_338, w_c4to2_carry_34_338, w_c4to2_cout_34_338;
math_compressor_4to2 u_c4to2_34_338 (
    .i_x1(w_c4to2_sum_34_240), .i_x2(w_c4to2_carry_33_333),
    .i_x3(w_c4to2_cout_33_333), .i_x4(w_c4to2_carry_33_334),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_338), .ow_carry(w_c4to2_carry_34_338), .ow_cout(w_c4to2_cout_34_338)
);
wire w_c4to2_sum_35_339, w_c4to2_carry_35_339, w_c4to2_cout_35_339;
math_compressor_4to2 u_c4to2_35_339 (
    .i_x1(w_c4to2_cout_34_238), .i_x2(w_c4to2_carry_34_239),
    .i_x3(w_c4to2_cout_34_239), .i_x4(w_c4to2_carry_34_240),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_339), .ow_carry(w_c4to2_carry_35_339), .ow_cout(w_c4to2_cout_35_339)
);
wire w_c4to2_sum_35_340, w_c4to2_carry_35_340, w_c4to2_cout_35_340;
math_compressor_4to2 u_c4to2_35_340 (
    .i_x1(w_c4to2_cout_34_240), .i_x2(w_c4to2_sum_35_241),
    .i_x3(w_c4to2_sum_35_242), .i_x4(w_c4to2_sum_35_243),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_340), .ow_carry(w_c4to2_carry_35_340), .ow_cout(w_c4to2_cout_35_340)
);
wire w_c4to2_sum_35_341, w_c4to2_carry_35_341, w_c4to2_cout_35_341;
math_compressor_4to2 u_c4to2_35_341 (
    .i_x1(w_c4to2_sum_35_244), .i_x2(w_c4to2_carry_34_336),
    .i_x3(w_c4to2_cout_34_336), .i_x4(w_c4to2_carry_34_337),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_341), .ow_carry(w_c4to2_carry_35_341), .ow_cout(w_c4to2_cout_35_341)
);
wire w_c4to2_sum_36_342, w_c4to2_carry_36_342, w_c4to2_cout_36_342;
math_compressor_4to2 u_c4to2_36_342 (
    .i_x1(w_c4to2_cout_35_242), .i_x2(w_c4to2_carry_35_243),
    .i_x3(w_c4to2_cout_35_243), .i_x4(w_c4to2_carry_35_244),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_342), .ow_carry(w_c4to2_carry_36_342), .ow_cout(w_c4to2_cout_36_342)
);
wire w_c4to2_sum_36_343, w_c4to2_carry_36_343, w_c4to2_cout_36_343;
math_compressor_4to2 u_c4to2_36_343 (
    .i_x1(w_c4to2_cout_35_244), .i_x2(w_c4to2_sum_36_245),
    .i_x3(w_c4to2_sum_36_246), .i_x4(w_c4to2_sum_36_247),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_343), .ow_carry(w_c4to2_carry_36_343), .ow_cout(w_c4to2_cout_36_343)
);
wire w_c4to2_sum_36_344, w_c4to2_carry_36_344, w_c4to2_cout_36_344;
math_compressor_4to2 u_c4to2_36_344 (
    .i_x1(w_c4to2_sum_36_248), .i_x2(w_c4to2_carry_35_339),
    .i_x3(w_c4to2_cout_35_339), .i_x4(w_c4to2_carry_35_340),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_344), .ow_carry(w_c4to2_carry_36_344), .ow_cout(w_c4to2_cout_36_344)
);
wire w_c4to2_sum_37_345, w_c4to2_carry_37_345, w_c4to2_cout_37_345;
math_compressor_4to2 u_c4to2_37_345 (
    .i_x1(w_c4to2_carry_36_246), .i_x2(w_c4to2_cout_36_246),
    .i_x3(w_c4to2_carry_36_247), .i_x4(w_c4to2_cout_36_247),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_345), .ow_carry(w_c4to2_carry_37_345), .ow_cout(w_c4to2_cout_37_345)
);
wire w_c4to2_sum_37_346, w_c4to2_carry_37_346, w_c4to2_cout_37_346;
math_compressor_4to2 u_c4to2_37_346 (
    .i_x1(w_c4to2_carry_36_248), .i_x2(w_c4to2_cout_36_248),
    .i_x3(w_c4to2_sum_37_249), .i_x4(w_c4to2_sum_37_250),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_346), .ow_carry(w_c4to2_carry_37_346), .ow_cout(w_c4to2_cout_37_346)
);
wire w_c4to2_sum_37_347, w_c4to2_carry_37_347, w_c4to2_cout_37_347;
math_compressor_4to2 u_c4to2_37_347 (
    .i_x1(w_c4to2_sum_37_251), .i_x2(w_c4to2_carry_36_342),
    .i_x3(w_c4to2_cout_36_342), .i_x4(w_c4to2_carry_36_343),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_347), .ow_carry(w_c4to2_carry_37_347), .ow_cout(w_c4to2_cout_37_347)
);
wire w_c4to2_sum_38_348, w_c4to2_carry_38_348, w_c4to2_cout_38_348;
math_compressor_4to2 u_c4to2_38_348 (
    .i_x1(w_pp_23_15), .i_x2(w_c4to2_carry_37_249),
    .i_x3(w_c4to2_cout_37_249), .i_x4(w_c4to2_carry_37_250),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_348), .ow_carry(w_c4to2_carry_38_348), .ow_cout(w_c4to2_cout_38_348)
);
wire w_c4to2_sum_38_349, w_c4to2_carry_38_349, w_c4to2_cout_38_349;
math_compressor_4to2 u_c4to2_38_349 (
    .i_x1(w_c4to2_cout_37_250), .i_x2(w_c4to2_carry_37_251),
    .i_x3(w_c4to2_cout_37_251), .i_x4(w_c4to2_sum_38_252),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_349), .ow_carry(w_c4to2_carry_38_349), .ow_cout(w_c4to2_cout_38_349)
);
wire w_c4to2_sum_38_350, w_c4to2_carry_38_350, w_c4to2_cout_38_350;
math_compressor_4to2 u_c4to2_38_350 (
    .i_x1(w_c4to2_sum_38_253), .i_x2(w_c4to2_carry_37_345),
    .i_x3(w_c4to2_cout_37_345), .i_x4(w_c4to2_carry_37_346),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_350), .ow_carry(w_c4to2_carry_38_350), .ow_cout(w_c4to2_cout_38_350)
);
wire w_c4to2_sum_39_351, w_c4to2_carry_39_351, w_c4to2_cout_39_351;
math_compressor_4to2 u_c4to2_39_351 (
    .i_x1(w_pp_20_19), .i_x2(w_pp_21_18),
    .i_x3(w_pp_22_17), .i_x4(w_pp_23_16),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_351), .ow_carry(w_c4to2_carry_39_351), .ow_cout(w_c4to2_cout_39_351)
);
wire w_c4to2_sum_39_352, w_c4to2_carry_39_352, w_c4to2_cout_39_352;
math_compressor_4to2 u_c4to2_39_352 (
    .i_x1(w_c4to2_carry_38_252), .i_x2(w_c4to2_cout_38_252),
    .i_x3(w_c4to2_carry_38_253), .i_x4(w_c4to2_cout_38_253),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_352), .ow_carry(w_c4to2_carry_39_352), .ow_cout(w_c4to2_cout_39_352)
);
wire w_c4to2_sum_39_353, w_c4to2_carry_39_353, w_c4to2_cout_39_353;
math_compressor_4to2 u_c4to2_39_353 (
    .i_x1(w_c4to2_sum_39_254), .i_x2(w_c4to2_carry_38_348),
    .i_x3(w_c4to2_cout_38_348), .i_x4(w_c4to2_carry_38_349),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_353), .ow_carry(w_c4to2_carry_39_353), .ow_cout(w_c4to2_cout_39_353)
);
wire w_c4to2_sum_40_354, w_c4to2_carry_40_354, w_c4to2_cout_40_354;
math_compressor_4to2 u_c4to2_40_354 (
    .i_x1(w_pp_17_23), .i_x2(w_pp_18_22),
    .i_x3(w_pp_19_21), .i_x4(w_pp_20_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_354), .ow_carry(w_c4to2_carry_40_354), .ow_cout(w_c4to2_cout_40_354)
);
wire w_c4to2_sum_40_355, w_c4to2_carry_40_355, w_c4to2_cout_40_355;
math_compressor_4to2 u_c4to2_40_355 (
    .i_x1(w_pp_21_19), .i_x2(w_pp_22_18),
    .i_x3(w_pp_23_17), .i_x4(w_c4to2_carry_39_254),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_355), .ow_carry(w_c4to2_carry_40_355), .ow_cout(w_c4to2_cout_40_355)
);
wire w_c4to2_sum_40_356, w_c4to2_carry_40_356, w_c4to2_cout_40_356;
math_compressor_4to2 u_c4to2_40_356 (
    .i_x1(w_c4to2_cout_39_254), .i_x2(w_c4to2_carry_39_351),
    .i_x3(w_c4to2_cout_39_351), .i_x4(w_c4to2_carry_39_352),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_356), .ow_carry(w_c4to2_carry_40_356), .ow_cout(w_c4to2_cout_40_356)
);
wire w_c4to2_sum_41_357, w_c4to2_carry_41_357, w_c4to2_cout_41_357;
math_compressor_4to2 u_c4to2_41_357 (
    .i_x1(w_pp_18_23), .i_x2(w_pp_19_22),
    .i_x3(w_pp_20_21), .i_x4(w_pp_21_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_357), .ow_carry(w_c4to2_carry_41_357), .ow_cout(w_c4to2_cout_41_357)
);
wire w_c4to2_sum_41_358, w_c4to2_carry_41_358, w_c4to2_cout_41_358;
math_compressor_4to2 u_c4to2_41_358 (
    .i_x1(w_pp_22_19), .i_x2(w_pp_23_18),
    .i_x3(w_c4to2_carry_40_354), .i_x4(w_c4to2_cout_40_354),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_358), .ow_carry(w_c4to2_carry_41_358), .ow_cout(w_c4to2_cout_41_358)
);
wire w_c4to2_sum_42_359, w_c4to2_carry_42_359, w_c4to2_cout_42_359;
math_compressor_4to2 u_c4to2_42_359 (
    .i_x1(w_pp_19_23), .i_x2(w_pp_20_22),
    .i_x3(w_pp_21_21), .i_x4(w_pp_22_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_42_359), .ow_carry(w_c4to2_carry_42_359), .ow_cout(w_c4to2_cout_42_359)
);

// Dadda Reduction Stage 5: height 6 -> 4

wire w_c4to2_sum_04_360, w_c4to2_carry_04_360, w_c4to2_cout_04_360;
math_compressor_4to2 u_c4to2_04_360 (
    .i_x1(w_pp_00_04), .i_x2(w_pp_01_03),
    .i_x3(w_pp_02_02), .i_x4(w_pp_03_01),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_04_360), .ow_carry(w_c4to2_carry_04_360), .ow_cout(w_c4to2_cout_04_360)
);
wire w_c4to2_sum_05_361, w_c4to2_carry_05_361, w_c4to2_cout_05_361;
math_compressor_4to2 u_c4to2_05_361 (
    .i_x1(w_pp_00_05), .i_x2(w_pp_01_04),
    .i_x3(w_pp_02_03), .i_x4(w_pp_03_02),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_05_361), .ow_carry(w_c4to2_carry_05_361), .ow_cout(w_c4to2_cout_05_361)
);
wire w_c4to2_sum_05_362, w_c4to2_carry_05_362, w_c4to2_cout_05_362;
math_compressor_4to2 u_c4to2_05_362 (
    .i_x1(w_pp_04_01), .i_x2(w_pp_05_00),
    .i_x3(w_c4to2_carry_04_360), .i_x4(w_c4to2_cout_04_360),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_05_362), .ow_carry(w_c4to2_carry_05_362), .ow_cout(w_c4to2_cout_05_362)
);
wire w_c4to2_sum_06_363, w_c4to2_carry_06_363, w_c4to2_cout_06_363;
math_compressor_4to2 u_c4to2_06_363 (
    .i_x1(w_pp_04_02), .i_x2(w_pp_05_01),
    .i_x3(w_pp_06_00), .i_x4(w_c4to2_sum_06_255),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_06_363), .ow_carry(w_c4to2_carry_06_363), .ow_cout(w_c4to2_cout_06_363)
);
wire w_c4to2_sum_06_364, w_c4to2_carry_06_364, w_c4to2_cout_06_364;
math_compressor_4to2 u_c4to2_06_364 (
    .i_x1(w_c4to2_carry_05_361), .i_x2(w_c4to2_cout_05_361),
    .i_x3(w_c4to2_carry_05_362), .i_x4(w_c4to2_cout_05_362),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_06_364), .ow_carry(w_c4to2_carry_06_364), .ow_cout(w_c4to2_cout_06_364)
);
wire w_c4to2_sum_07_365, w_c4to2_carry_07_365, w_c4to2_cout_07_365;
math_compressor_4to2 u_c4to2_07_365 (
    .i_x1(w_c4to2_carry_06_255), .i_x2(w_c4to2_cout_06_255),
    .i_x3(w_c4to2_sum_07_256), .i_x4(w_c4to2_sum_07_257),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_07_365), .ow_carry(w_c4to2_carry_07_365), .ow_cout(w_c4to2_cout_07_365)
);
wire w_c4to2_sum_07_366, w_c4to2_carry_07_366, w_c4to2_cout_07_366;
math_compressor_4to2 u_c4to2_07_366 (
    .i_x1(w_c4to2_carry_06_363), .i_x2(w_c4to2_cout_06_363),
    .i_x3(w_c4to2_carry_06_364), .i_x4(w_c4to2_cout_06_364),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_07_366), .ow_carry(w_c4to2_carry_07_366), .ow_cout(w_c4to2_cout_07_366)
);
wire w_c4to2_sum_08_367, w_c4to2_carry_08_367, w_c4to2_cout_08_367;
math_compressor_4to2 u_c4to2_08_367 (
    .i_x1(w_c4to2_cout_07_257), .i_x2(w_c4to2_sum_08_258),
    .i_x3(w_c4to2_sum_08_259), .i_x4(w_c4to2_sum_08_260),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_367), .ow_carry(w_c4to2_carry_08_367), .ow_cout(w_c4to2_cout_08_367)
);
wire w_c4to2_sum_08_368, w_c4to2_carry_08_368, w_c4to2_cout_08_368;
math_compressor_4to2 u_c4to2_08_368 (
    .i_x1(w_c4to2_carry_07_365), .i_x2(w_c4to2_cout_07_365),
    .i_x3(w_c4to2_carry_07_366), .i_x4(w_c4to2_cout_07_366),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_368), .ow_carry(w_c4to2_carry_08_368), .ow_cout(w_c4to2_cout_08_368)
);
wire w_c4to2_sum_09_369, w_c4to2_carry_09_369, w_c4to2_cout_09_369;
math_compressor_4to2 u_c4to2_09_369 (
    .i_x1(w_c4to2_cout_08_260), .i_x2(w_c4to2_sum_09_261),
    .i_x3(w_c4to2_sum_09_262), .i_x4(w_c4to2_sum_09_263),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_369), .ow_carry(w_c4to2_carry_09_369), .ow_cout(w_c4to2_cout_09_369)
);
wire w_c4to2_sum_09_370, w_c4to2_carry_09_370, w_c4to2_cout_09_370;
math_compressor_4to2 u_c4to2_09_370 (
    .i_x1(w_c4to2_carry_08_367), .i_x2(w_c4to2_cout_08_367),
    .i_x3(w_c4to2_carry_08_368), .i_x4(w_c4to2_cout_08_368),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_370), .ow_carry(w_c4to2_carry_09_370), .ow_cout(w_c4to2_cout_09_370)
);
wire w_c4to2_sum_10_371, w_c4to2_carry_10_371, w_c4to2_cout_10_371;
math_compressor_4to2 u_c4to2_10_371 (
    .i_x1(w_c4to2_cout_09_263), .i_x2(w_c4to2_sum_10_264),
    .i_x3(w_c4to2_sum_10_265), .i_x4(w_c4to2_sum_10_266),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_371), .ow_carry(w_c4to2_carry_10_371), .ow_cout(w_c4to2_cout_10_371)
);
wire w_c4to2_sum_10_372, w_c4to2_carry_10_372, w_c4to2_cout_10_372;
math_compressor_4to2 u_c4to2_10_372 (
    .i_x1(w_c4to2_carry_09_369), .i_x2(w_c4to2_cout_09_369),
    .i_x3(w_c4to2_carry_09_370), .i_x4(w_c4to2_cout_09_370),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_372), .ow_carry(w_c4to2_carry_10_372), .ow_cout(w_c4to2_cout_10_372)
);
wire w_c4to2_sum_11_373, w_c4to2_carry_11_373, w_c4to2_cout_11_373;
math_compressor_4to2 u_c4to2_11_373 (
    .i_x1(w_c4to2_cout_10_266), .i_x2(w_c4to2_sum_11_267),
    .i_x3(w_c4to2_sum_11_268), .i_x4(w_c4to2_sum_11_269),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_373), .ow_carry(w_c4to2_carry_11_373), .ow_cout(w_c4to2_cout_11_373)
);
wire w_c4to2_sum_11_374, w_c4to2_carry_11_374, w_c4to2_cout_11_374;
math_compressor_4to2 u_c4to2_11_374 (
    .i_x1(w_c4to2_carry_10_371), .i_x2(w_c4to2_cout_10_371),
    .i_x3(w_c4to2_carry_10_372), .i_x4(w_c4to2_cout_10_372),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_374), .ow_carry(w_c4to2_carry_11_374), .ow_cout(w_c4to2_cout_11_374)
);
wire w_c4to2_sum_12_375, w_c4to2_carry_12_375, w_c4to2_cout_12_375;
math_compressor_4to2 u_c4to2_12_375 (
    .i_x1(w_c4to2_cout_11_269), .i_x2(w_c4to2_sum_12_270),
    .i_x3(w_c4to2_sum_12_271), .i_x4(w_c4to2_sum_12_272),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_375), .ow_carry(w_c4to2_carry_12_375), .ow_cout(w_c4to2_cout_12_375)
);
wire w_c4to2_sum_12_376, w_c4to2_carry_12_376, w_c4to2_cout_12_376;
math_compressor_4to2 u_c4to2_12_376 (
    .i_x1(w_c4to2_carry_11_373), .i_x2(w_c4to2_cout_11_373),
    .i_x3(w_c4to2_carry_11_374), .i_x4(w_c4to2_cout_11_374),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_376), .ow_carry(w_c4to2_carry_12_376), .ow_cout(w_c4to2_cout_12_376)
);
wire w_c4to2_sum_13_377, w_c4to2_carry_13_377, w_c4to2_cout_13_377;
math_compressor_4to2 u_c4to2_13_377 (
    .i_x1(w_c4to2_cout_12_272), .i_x2(w_c4to2_sum_13_273),
    .i_x3(w_c4to2_sum_13_274), .i_x4(w_c4to2_sum_13_275),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_377), .ow_carry(w_c4to2_carry_13_377), .ow_cout(w_c4to2_cout_13_377)
);
wire w_c4to2_sum_13_378, w_c4to2_carry_13_378, w_c4to2_cout_13_378;
math_compressor_4to2 u_c4to2_13_378 (
    .i_x1(w_c4to2_carry_12_375), .i_x2(w_c4to2_cout_12_375),
    .i_x3(w_c4to2_carry_12_376), .i_x4(w_c4to2_cout_12_376),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_378), .ow_carry(w_c4to2_carry_13_378), .ow_cout(w_c4to2_cout_13_378)
);
wire w_c4to2_sum_14_379, w_c4to2_carry_14_379, w_c4to2_cout_14_379;
math_compressor_4to2 u_c4to2_14_379 (
    .i_x1(w_c4to2_cout_13_275), .i_x2(w_c4to2_sum_14_276),
    .i_x3(w_c4to2_sum_14_277), .i_x4(w_c4to2_sum_14_278),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_379), .ow_carry(w_c4to2_carry_14_379), .ow_cout(w_c4to2_cout_14_379)
);
wire w_c4to2_sum_14_380, w_c4to2_carry_14_380, w_c4to2_cout_14_380;
math_compressor_4to2 u_c4to2_14_380 (
    .i_x1(w_c4to2_carry_13_377), .i_x2(w_c4to2_cout_13_377),
    .i_x3(w_c4to2_carry_13_378), .i_x4(w_c4to2_cout_13_378),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_380), .ow_carry(w_c4to2_carry_14_380), .ow_cout(w_c4to2_cout_14_380)
);
wire w_c4to2_sum_15_381, w_c4to2_carry_15_381, w_c4to2_cout_15_381;
math_compressor_4to2 u_c4to2_15_381 (
    .i_x1(w_c4to2_cout_14_278), .i_x2(w_c4to2_sum_15_279),
    .i_x3(w_c4to2_sum_15_280), .i_x4(w_c4to2_sum_15_281),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_381), .ow_carry(w_c4to2_carry_15_381), .ow_cout(w_c4to2_cout_15_381)
);
wire w_c4to2_sum_15_382, w_c4to2_carry_15_382, w_c4to2_cout_15_382;
math_compressor_4to2 u_c4to2_15_382 (
    .i_x1(w_c4to2_carry_14_379), .i_x2(w_c4to2_cout_14_379),
    .i_x3(w_c4to2_carry_14_380), .i_x4(w_c4to2_cout_14_380),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_382), .ow_carry(w_c4to2_carry_15_382), .ow_cout(w_c4to2_cout_15_382)
);
wire w_c4to2_sum_16_383, w_c4to2_carry_16_383, w_c4to2_cout_16_383;
math_compressor_4to2 u_c4to2_16_383 (
    .i_x1(w_c4to2_cout_15_281), .i_x2(w_c4to2_sum_16_282),
    .i_x3(w_c4to2_sum_16_283), .i_x4(w_c4to2_sum_16_284),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_383), .ow_carry(w_c4to2_carry_16_383), .ow_cout(w_c4to2_cout_16_383)
);
wire w_c4to2_sum_16_384, w_c4to2_carry_16_384, w_c4to2_cout_16_384;
math_compressor_4to2 u_c4to2_16_384 (
    .i_x1(w_c4to2_carry_15_381), .i_x2(w_c4to2_cout_15_381),
    .i_x3(w_c4to2_carry_15_382), .i_x4(w_c4to2_cout_15_382),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_384), .ow_carry(w_c4to2_carry_16_384), .ow_cout(w_c4to2_cout_16_384)
);
wire w_c4to2_sum_17_385, w_c4to2_carry_17_385, w_c4to2_cout_17_385;
math_compressor_4to2 u_c4to2_17_385 (
    .i_x1(w_c4to2_cout_16_284), .i_x2(w_c4to2_sum_17_285),
    .i_x3(w_c4to2_sum_17_286), .i_x4(w_c4to2_sum_17_287),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_385), .ow_carry(w_c4to2_carry_17_385), .ow_cout(w_c4to2_cout_17_385)
);
wire w_c4to2_sum_17_386, w_c4to2_carry_17_386, w_c4to2_cout_17_386;
math_compressor_4to2 u_c4to2_17_386 (
    .i_x1(w_c4to2_carry_16_383), .i_x2(w_c4to2_cout_16_383),
    .i_x3(w_c4to2_carry_16_384), .i_x4(w_c4to2_cout_16_384),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_386), .ow_carry(w_c4to2_carry_17_386), .ow_cout(w_c4to2_cout_17_386)
);
wire w_c4to2_sum_18_387, w_c4to2_carry_18_387, w_c4to2_cout_18_387;
math_compressor_4to2 u_c4to2_18_387 (
    .i_x1(w_c4to2_cout_17_287), .i_x2(w_c4to2_sum_18_288),
    .i_x3(w_c4to2_sum_18_289), .i_x4(w_c4to2_sum_18_290),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_387), .ow_carry(w_c4to2_carry_18_387), .ow_cout(w_c4to2_cout_18_387)
);
wire w_c4to2_sum_18_388, w_c4to2_carry_18_388, w_c4to2_cout_18_388;
math_compressor_4to2 u_c4to2_18_388 (
    .i_x1(w_c4to2_carry_17_385), .i_x2(w_c4to2_cout_17_385),
    .i_x3(w_c4to2_carry_17_386), .i_x4(w_c4to2_cout_17_386),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_388), .ow_carry(w_c4to2_carry_18_388), .ow_cout(w_c4to2_cout_18_388)
);
wire w_c4to2_sum_19_389, w_c4to2_carry_19_389, w_c4to2_cout_19_389;
math_compressor_4to2 u_c4to2_19_389 (
    .i_x1(w_c4to2_cout_18_290), .i_x2(w_c4to2_sum_19_291),
    .i_x3(w_c4to2_sum_19_292), .i_x4(w_c4to2_sum_19_293),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_389), .ow_carry(w_c4to2_carry_19_389), .ow_cout(w_c4to2_cout_19_389)
);
wire w_c4to2_sum_19_390, w_c4to2_carry_19_390, w_c4to2_cout_19_390;
math_compressor_4to2 u_c4to2_19_390 (
    .i_x1(w_c4to2_carry_18_387), .i_x2(w_c4to2_cout_18_387),
    .i_x3(w_c4to2_carry_18_388), .i_x4(w_c4to2_cout_18_388),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_390), .ow_carry(w_c4to2_carry_19_390), .ow_cout(w_c4to2_cout_19_390)
);
wire w_c4to2_sum_20_391, w_c4to2_carry_20_391, w_c4to2_cout_20_391;
math_compressor_4to2 u_c4to2_20_391 (
    .i_x1(w_c4to2_cout_19_293), .i_x2(w_c4to2_sum_20_294),
    .i_x3(w_c4to2_sum_20_295), .i_x4(w_c4to2_sum_20_296),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_391), .ow_carry(w_c4to2_carry_20_391), .ow_cout(w_c4to2_cout_20_391)
);
wire w_c4to2_sum_20_392, w_c4to2_carry_20_392, w_c4to2_cout_20_392;
math_compressor_4to2 u_c4to2_20_392 (
    .i_x1(w_c4to2_carry_19_389), .i_x2(w_c4to2_cout_19_389),
    .i_x3(w_c4to2_carry_19_390), .i_x4(w_c4to2_cout_19_390),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_392), .ow_carry(w_c4to2_carry_20_392), .ow_cout(w_c4to2_cout_20_392)
);
wire w_c4to2_sum_21_393, w_c4to2_carry_21_393, w_c4to2_cout_21_393;
math_compressor_4to2 u_c4to2_21_393 (
    .i_x1(w_c4to2_cout_20_296), .i_x2(w_c4to2_sum_21_297),
    .i_x3(w_c4to2_sum_21_298), .i_x4(w_c4to2_sum_21_299),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_393), .ow_carry(w_c4to2_carry_21_393), .ow_cout(w_c4to2_cout_21_393)
);
wire w_c4to2_sum_21_394, w_c4to2_carry_21_394, w_c4to2_cout_21_394;
math_compressor_4to2 u_c4to2_21_394 (
    .i_x1(w_c4to2_carry_20_391), .i_x2(w_c4to2_cout_20_391),
    .i_x3(w_c4to2_carry_20_392), .i_x4(w_c4to2_cout_20_392),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_394), .ow_carry(w_c4to2_carry_21_394), .ow_cout(w_c4to2_cout_21_394)
);
wire w_c4to2_sum_22_395, w_c4to2_carry_22_395, w_c4to2_cout_22_395;
math_compressor_4to2 u_c4to2_22_395 (
    .i_x1(w_c4to2_cout_21_299), .i_x2(w_c4to2_sum_22_300),
    .i_x3(w_c4to2_sum_22_301), .i_x4(w_c4to2_sum_22_302),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_395), .ow_carry(w_c4to2_carry_22_395), .ow_cout(w_c4to2_cout_22_395)
);
wire w_c4to2_sum_22_396, w_c4to2_carry_22_396, w_c4to2_cout_22_396;
math_compressor_4to2 u_c4to2_22_396 (
    .i_x1(w_c4to2_carry_21_393), .i_x2(w_c4to2_cout_21_393),
    .i_x3(w_c4to2_carry_21_394), .i_x4(w_c4to2_cout_21_394),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_396), .ow_carry(w_c4to2_carry_22_396), .ow_cout(w_c4to2_cout_22_396)
);
wire w_c4to2_sum_23_397, w_c4to2_carry_23_397, w_c4to2_cout_23_397;
math_compressor_4to2 u_c4to2_23_397 (
    .i_x1(w_c4to2_cout_22_302), .i_x2(w_c4to2_sum_23_303),
    .i_x3(w_c4to2_sum_23_304), .i_x4(w_c4to2_sum_23_305),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_397), .ow_carry(w_c4to2_carry_23_397), .ow_cout(w_c4to2_cout_23_397)
);
wire w_c4to2_sum_23_398, w_c4to2_carry_23_398, w_c4to2_cout_23_398;
math_compressor_4to2 u_c4to2_23_398 (
    .i_x1(w_c4to2_carry_22_395), .i_x2(w_c4to2_cout_22_395),
    .i_x3(w_c4to2_carry_22_396), .i_x4(w_c4to2_cout_22_396),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_398), .ow_carry(w_c4to2_carry_23_398), .ow_cout(w_c4to2_cout_23_398)
);
wire w_c4to2_sum_24_399, w_c4to2_carry_24_399, w_c4to2_cout_24_399;
math_compressor_4to2 u_c4to2_24_399 (
    .i_x1(w_c4to2_carry_23_305), .i_x2(w_c4to2_cout_23_305),
    .i_x3(w_c4to2_sum_24_306), .i_x4(w_c4to2_sum_24_307),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_399), .ow_carry(w_c4to2_carry_24_399), .ow_cout(w_c4to2_cout_24_399)
);
wire w_c4to2_sum_24_400, w_c4to2_carry_24_400, w_c4to2_cout_24_400;
math_compressor_4to2 u_c4to2_24_400 (
    .i_x1(w_c4to2_sum_24_308), .i_x2(w_c4to2_carry_23_397),
    .i_x3(w_c4to2_cout_23_397), .i_x4(w_c4to2_carry_23_398),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_400), .ow_carry(w_c4to2_carry_24_400), .ow_cout(w_c4to2_cout_24_400)
);
wire w_c4to2_sum_25_401, w_c4to2_carry_25_401, w_c4to2_cout_25_401;
math_compressor_4to2 u_c4to2_25_401 (
    .i_x1(w_c4to2_cout_24_308), .i_x2(w_c4to2_sum_25_309),
    .i_x3(w_c4to2_sum_25_310), .i_x4(w_c4to2_sum_25_311),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_401), .ow_carry(w_c4to2_carry_25_401), .ow_cout(w_c4to2_cout_25_401)
);
wire w_c4to2_sum_25_402, w_c4to2_carry_25_402, w_c4to2_cout_25_402;
math_compressor_4to2 u_c4to2_25_402 (
    .i_x1(w_c4to2_carry_24_399), .i_x2(w_c4to2_cout_24_399),
    .i_x3(w_c4to2_carry_24_400), .i_x4(w_c4to2_cout_24_400),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_402), .ow_carry(w_c4to2_carry_25_402), .ow_cout(w_c4to2_cout_25_402)
);
wire w_c4to2_sum_26_403, w_c4to2_carry_26_403, w_c4to2_cout_26_403;
math_compressor_4to2 u_c4to2_26_403 (
    .i_x1(w_c4to2_cout_25_310), .i_x2(w_c4to2_carry_25_311),
    .i_x3(w_c4to2_cout_25_311), .i_x4(w_c4to2_sum_26_312),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_403), .ow_carry(w_c4to2_carry_26_403), .ow_cout(w_c4to2_cout_26_403)
);
wire w_c4to2_sum_26_404, w_c4to2_carry_26_404, w_c4to2_cout_26_404;
math_compressor_4to2 u_c4to2_26_404 (
    .i_x1(w_c4to2_sum_26_313), .i_x2(w_c4to2_sum_26_314),
    .i_x3(w_c4to2_carry_25_401), .i_x4(w_c4to2_cout_25_401),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_404), .ow_carry(w_c4to2_carry_26_404), .ow_cout(w_c4to2_cout_26_404)
);
wire w_c4to2_sum_27_405, w_c4to2_carry_27_405, w_c4to2_cout_27_405;
math_compressor_4to2 u_c4to2_27_405 (
    .i_x1(w_c4to2_cout_26_313), .i_x2(w_c4to2_carry_26_314),
    .i_x3(w_c4to2_cout_26_314), .i_x4(w_c4to2_sum_27_315),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_405), .ow_carry(w_c4to2_carry_27_405), .ow_cout(w_c4to2_cout_27_405)
);
wire w_c4to2_sum_27_406, w_c4to2_carry_27_406, w_c4to2_cout_27_406;
math_compressor_4to2 u_c4to2_27_406 (
    .i_x1(w_c4to2_sum_27_316), .i_x2(w_c4to2_sum_27_317),
    .i_x3(w_c4to2_carry_26_403), .i_x4(w_c4to2_cout_26_403),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_406), .ow_carry(w_c4to2_carry_27_406), .ow_cout(w_c4to2_cout_27_406)
);
wire w_c4to2_sum_28_407, w_c4to2_carry_28_407, w_c4to2_cout_28_407;
math_compressor_4to2 u_c4to2_28_407 (
    .i_x1(w_c4to2_cout_27_316), .i_x2(w_c4to2_carry_27_317),
    .i_x3(w_c4to2_cout_27_317), .i_x4(w_c4to2_sum_28_318),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_407), .ow_carry(w_c4to2_carry_28_407), .ow_cout(w_c4to2_cout_28_407)
);
wire w_c4to2_sum_28_408, w_c4to2_carry_28_408, w_c4to2_cout_28_408;
math_compressor_4to2 u_c4to2_28_408 (
    .i_x1(w_c4to2_sum_28_319), .i_x2(w_c4to2_sum_28_320),
    .i_x3(w_c4to2_carry_27_405), .i_x4(w_c4to2_cout_27_405),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_408), .ow_carry(w_c4to2_carry_28_408), .ow_cout(w_c4to2_cout_28_408)
);
wire w_c4to2_sum_29_409, w_c4to2_carry_29_409, w_c4to2_cout_29_409;
math_compressor_4to2 u_c4to2_29_409 (
    .i_x1(w_c4to2_cout_28_319), .i_x2(w_c4to2_carry_28_320),
    .i_x3(w_c4to2_cout_28_320), .i_x4(w_c4to2_sum_29_321),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_409), .ow_carry(w_c4to2_carry_29_409), .ow_cout(w_c4to2_cout_29_409)
);
wire w_c4to2_sum_29_410, w_c4to2_carry_29_410, w_c4to2_cout_29_410;
math_compressor_4to2 u_c4to2_29_410 (
    .i_x1(w_c4to2_sum_29_322), .i_x2(w_c4to2_sum_29_323),
    .i_x3(w_c4to2_carry_28_407), .i_x4(w_c4to2_cout_28_407),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_410), .ow_carry(w_c4to2_carry_29_410), .ow_cout(w_c4to2_cout_29_410)
);
wire w_c4to2_sum_30_411, w_c4to2_carry_30_411, w_c4to2_cout_30_411;
math_compressor_4to2 u_c4to2_30_411 (
    .i_x1(w_c4to2_cout_29_322), .i_x2(w_c4to2_carry_29_323),
    .i_x3(w_c4to2_cout_29_323), .i_x4(w_c4to2_sum_30_324),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_411), .ow_carry(w_c4to2_carry_30_411), .ow_cout(w_c4to2_cout_30_411)
);
wire w_c4to2_sum_30_412, w_c4to2_carry_30_412, w_c4to2_cout_30_412;
math_compressor_4to2 u_c4to2_30_412 (
    .i_x1(w_c4to2_sum_30_325), .i_x2(w_c4to2_sum_30_326),
    .i_x3(w_c4to2_carry_29_409), .i_x4(w_c4to2_cout_29_409),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_412), .ow_carry(w_c4to2_carry_30_412), .ow_cout(w_c4to2_cout_30_412)
);
wire w_c4to2_sum_31_413, w_c4to2_carry_31_413, w_c4to2_cout_31_413;
math_compressor_4to2 u_c4to2_31_413 (
    .i_x1(w_c4to2_cout_30_325), .i_x2(w_c4to2_carry_30_326),
    .i_x3(w_c4to2_cout_30_326), .i_x4(w_c4to2_sum_31_327),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_413), .ow_carry(w_c4to2_carry_31_413), .ow_cout(w_c4to2_cout_31_413)
);
wire w_c4to2_sum_31_414, w_c4to2_carry_31_414, w_c4to2_cout_31_414;
math_compressor_4to2 u_c4to2_31_414 (
    .i_x1(w_c4to2_sum_31_328), .i_x2(w_c4to2_sum_31_329),
    .i_x3(w_c4to2_carry_30_411), .i_x4(w_c4to2_cout_30_411),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_414), .ow_carry(w_c4to2_carry_31_414), .ow_cout(w_c4to2_cout_31_414)
);
wire w_c4to2_sum_32_415, w_c4to2_carry_32_415, w_c4to2_cout_32_415;
math_compressor_4to2 u_c4to2_32_415 (
    .i_x1(w_c4to2_cout_31_328), .i_x2(w_c4to2_carry_31_329),
    .i_x3(w_c4to2_cout_31_329), .i_x4(w_c4to2_sum_32_330),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_415), .ow_carry(w_c4to2_carry_32_415), .ow_cout(w_c4to2_cout_32_415)
);
wire w_c4to2_sum_32_416, w_c4to2_carry_32_416, w_c4to2_cout_32_416;
math_compressor_4to2 u_c4to2_32_416 (
    .i_x1(w_c4to2_sum_32_331), .i_x2(w_c4to2_sum_32_332),
    .i_x3(w_c4to2_carry_31_413), .i_x4(w_c4to2_cout_31_413),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_416), .ow_carry(w_c4to2_carry_32_416), .ow_cout(w_c4to2_cout_32_416)
);
wire w_c4to2_sum_33_417, w_c4to2_carry_33_417, w_c4to2_cout_33_417;
math_compressor_4to2 u_c4to2_33_417 (
    .i_x1(w_c4to2_cout_32_331), .i_x2(w_c4to2_carry_32_332),
    .i_x3(w_c4to2_cout_32_332), .i_x4(w_c4to2_sum_33_333),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_417), .ow_carry(w_c4to2_carry_33_417), .ow_cout(w_c4to2_cout_33_417)
);
wire w_c4to2_sum_33_418, w_c4to2_carry_33_418, w_c4to2_cout_33_418;
math_compressor_4to2 u_c4to2_33_418 (
    .i_x1(w_c4to2_sum_33_334), .i_x2(w_c4to2_sum_33_335),
    .i_x3(w_c4to2_carry_32_415), .i_x4(w_c4to2_cout_32_415),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_418), .ow_carry(w_c4to2_carry_33_418), .ow_cout(w_c4to2_cout_33_418)
);
wire w_c4to2_sum_34_419, w_c4to2_carry_34_419, w_c4to2_cout_34_419;
math_compressor_4to2 u_c4to2_34_419 (
    .i_x1(w_c4to2_cout_33_334), .i_x2(w_c4to2_carry_33_335),
    .i_x3(w_c4to2_cout_33_335), .i_x4(w_c4to2_sum_34_336),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_419), .ow_carry(w_c4to2_carry_34_419), .ow_cout(w_c4to2_cout_34_419)
);
wire w_c4to2_sum_34_420, w_c4to2_carry_34_420, w_c4to2_cout_34_420;
math_compressor_4to2 u_c4to2_34_420 (
    .i_x1(w_c4to2_sum_34_337), .i_x2(w_c4to2_sum_34_338),
    .i_x3(w_c4to2_carry_33_417), .i_x4(w_c4to2_cout_33_417),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_420), .ow_carry(w_c4to2_carry_34_420), .ow_cout(w_c4to2_cout_34_420)
);
wire w_c4to2_sum_35_421, w_c4to2_carry_35_421, w_c4to2_cout_35_421;
math_compressor_4to2 u_c4to2_35_421 (
    .i_x1(w_c4to2_cout_34_337), .i_x2(w_c4to2_carry_34_338),
    .i_x3(w_c4to2_cout_34_338), .i_x4(w_c4to2_sum_35_339),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_421), .ow_carry(w_c4to2_carry_35_421), .ow_cout(w_c4to2_cout_35_421)
);
wire w_c4to2_sum_35_422, w_c4to2_carry_35_422, w_c4to2_cout_35_422;
math_compressor_4to2 u_c4to2_35_422 (
    .i_x1(w_c4to2_sum_35_340), .i_x2(w_c4to2_sum_35_341),
    .i_x3(w_c4to2_carry_34_419), .i_x4(w_c4to2_cout_34_419),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_422), .ow_carry(w_c4to2_carry_35_422), .ow_cout(w_c4to2_cout_35_422)
);
wire w_c4to2_sum_36_423, w_c4to2_carry_36_423, w_c4to2_cout_36_423;
math_compressor_4to2 u_c4to2_36_423 (
    .i_x1(w_c4to2_cout_35_340), .i_x2(w_c4to2_carry_35_341),
    .i_x3(w_c4to2_cout_35_341), .i_x4(w_c4to2_sum_36_342),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_423), .ow_carry(w_c4to2_carry_36_423), .ow_cout(w_c4to2_cout_36_423)
);
wire w_c4to2_sum_36_424, w_c4to2_carry_36_424, w_c4to2_cout_36_424;
math_compressor_4to2 u_c4to2_36_424 (
    .i_x1(w_c4to2_sum_36_343), .i_x2(w_c4to2_sum_36_344),
    .i_x3(w_c4to2_carry_35_421), .i_x4(w_c4to2_cout_35_421),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_424), .ow_carry(w_c4to2_carry_36_424), .ow_cout(w_c4to2_cout_36_424)
);
wire w_c4to2_sum_37_425, w_c4to2_carry_37_425, w_c4to2_cout_37_425;
math_compressor_4to2 u_c4to2_37_425 (
    .i_x1(w_c4to2_cout_36_343), .i_x2(w_c4to2_carry_36_344),
    .i_x3(w_c4to2_cout_36_344), .i_x4(w_c4to2_sum_37_345),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_425), .ow_carry(w_c4to2_carry_37_425), .ow_cout(w_c4to2_cout_37_425)
);
wire w_c4to2_sum_37_426, w_c4to2_carry_37_426, w_c4to2_cout_37_426;
math_compressor_4to2 u_c4to2_37_426 (
    .i_x1(w_c4to2_sum_37_346), .i_x2(w_c4to2_sum_37_347),
    .i_x3(w_c4to2_carry_36_423), .i_x4(w_c4to2_cout_36_423),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_426), .ow_carry(w_c4to2_carry_37_426), .ow_cout(w_c4to2_cout_37_426)
);
wire w_c4to2_sum_38_427, w_c4to2_carry_38_427, w_c4to2_cout_38_427;
math_compressor_4to2 u_c4to2_38_427 (
    .i_x1(w_c4to2_cout_37_346), .i_x2(w_c4to2_carry_37_347),
    .i_x3(w_c4to2_cout_37_347), .i_x4(w_c4to2_sum_38_348),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_427), .ow_carry(w_c4to2_carry_38_427), .ow_cout(w_c4to2_cout_38_427)
);
wire w_c4to2_sum_38_428, w_c4to2_carry_38_428, w_c4to2_cout_38_428;
math_compressor_4to2 u_c4to2_38_428 (
    .i_x1(w_c4to2_sum_38_349), .i_x2(w_c4to2_sum_38_350),
    .i_x3(w_c4to2_carry_37_425), .i_x4(w_c4to2_cout_37_425),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_428), .ow_carry(w_c4to2_carry_38_428), .ow_cout(w_c4to2_cout_38_428)
);
wire w_c4to2_sum_39_429, w_c4to2_carry_39_429, w_c4to2_cout_39_429;
math_compressor_4to2 u_c4to2_39_429 (
    .i_x1(w_c4to2_cout_38_349), .i_x2(w_c4to2_carry_38_350),
    .i_x3(w_c4to2_cout_38_350), .i_x4(w_c4to2_sum_39_351),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_429), .ow_carry(w_c4to2_carry_39_429), .ow_cout(w_c4to2_cout_39_429)
);
wire w_c4to2_sum_39_430, w_c4to2_carry_39_430, w_c4to2_cout_39_430;
math_compressor_4to2 u_c4to2_39_430 (
    .i_x1(w_c4to2_sum_39_352), .i_x2(w_c4to2_sum_39_353),
    .i_x3(w_c4to2_carry_38_427), .i_x4(w_c4to2_cout_38_427),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_430), .ow_carry(w_c4to2_carry_39_430), .ow_cout(w_c4to2_cout_39_430)
);
wire w_c4to2_sum_40_431, w_c4to2_carry_40_431, w_c4to2_cout_40_431;
math_compressor_4to2 u_c4to2_40_431 (
    .i_x1(w_c4to2_cout_39_352), .i_x2(w_c4to2_carry_39_353),
    .i_x3(w_c4to2_cout_39_353), .i_x4(w_c4to2_sum_40_354),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_431), .ow_carry(w_c4to2_carry_40_431), .ow_cout(w_c4to2_cout_40_431)
);
wire w_c4to2_sum_40_432, w_c4to2_carry_40_432, w_c4to2_cout_40_432;
math_compressor_4to2 u_c4to2_40_432 (
    .i_x1(w_c4to2_sum_40_355), .i_x2(w_c4to2_sum_40_356),
    .i_x3(w_c4to2_carry_39_429), .i_x4(w_c4to2_cout_39_429),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_432), .ow_carry(w_c4to2_carry_40_432), .ow_cout(w_c4to2_cout_40_432)
);
wire w_c4to2_sum_41_433, w_c4to2_carry_41_433, w_c4to2_cout_41_433;
math_compressor_4to2 u_c4to2_41_433 (
    .i_x1(w_c4to2_carry_40_355), .i_x2(w_c4to2_cout_40_355),
    .i_x3(w_c4to2_carry_40_356), .i_x4(w_c4to2_cout_40_356),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_433), .ow_carry(w_c4to2_carry_41_433), .ow_cout(w_c4to2_cout_41_433)
);
wire w_c4to2_sum_41_434, w_c4to2_carry_41_434, w_c4to2_cout_41_434;
math_compressor_4to2 u_c4to2_41_434 (
    .i_x1(w_c4to2_sum_41_357), .i_x2(w_c4to2_sum_41_358),
    .i_x3(w_c4to2_carry_40_431), .i_x4(w_c4to2_cout_40_431),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_434), .ow_carry(w_c4to2_carry_41_434), .ow_cout(w_c4to2_cout_41_434)
);
wire w_c4to2_sum_42_435, w_c4to2_carry_42_435, w_c4to2_cout_42_435;
math_compressor_4to2 u_c4to2_42_435 (
    .i_x1(w_pp_23_19), .i_x2(w_c4to2_carry_41_357),
    .i_x3(w_c4to2_cout_41_357), .i_x4(w_c4to2_carry_41_358),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_42_435), .ow_carry(w_c4to2_carry_42_435), .ow_cout(w_c4to2_cout_42_435)
);
wire w_c4to2_sum_42_436, w_c4to2_carry_42_436, w_c4to2_cout_42_436;
math_compressor_4to2 u_c4to2_42_436 (
    .i_x1(w_c4to2_cout_41_358), .i_x2(w_c4to2_sum_42_359),
    .i_x3(w_c4to2_carry_41_433), .i_x4(w_c4to2_cout_41_433),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_42_436), .ow_carry(w_c4to2_carry_42_436), .ow_cout(w_c4to2_cout_42_436)
);
wire w_c4to2_sum_43_437, w_c4to2_carry_43_437, w_c4to2_cout_43_437;
math_compressor_4to2 u_c4to2_43_437 (
    .i_x1(w_pp_20_23), .i_x2(w_pp_21_22),
    .i_x3(w_pp_22_21), .i_x4(w_pp_23_20),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_43_437), .ow_carry(w_c4to2_carry_43_437), .ow_cout(w_c4to2_cout_43_437)
);
wire w_c4to2_sum_43_438, w_c4to2_carry_43_438, w_c4to2_cout_43_438;
math_compressor_4to2 u_c4to2_43_438 (
    .i_x1(w_c4to2_carry_42_359), .i_x2(w_c4to2_cout_42_359),
    .i_x3(w_c4to2_carry_42_435), .i_x4(w_c4to2_cout_42_435),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_43_438), .ow_carry(w_c4to2_carry_43_438), .ow_cout(w_c4to2_cout_43_438)
);
wire w_c4to2_sum_44_439, w_c4to2_carry_44_439, w_c4to2_cout_44_439;
math_compressor_4to2 u_c4to2_44_439 (
    .i_x1(w_pp_21_23), .i_x2(w_pp_22_22),
    .i_x3(w_pp_23_21), .i_x4(w_c4to2_carry_43_437),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_44_439), .ow_carry(w_c4to2_carry_44_439), .ow_cout(w_c4to2_cout_44_439)
);

// Dadda Reduction Stage 6: height 4 -> 3

wire w_c4to2_sum_03_440, w_c4to2_carry_03_440, w_c4to2_cout_03_440;
math_compressor_4to2 u_c4to2_03_440 (
    .i_x1(w_pp_00_03), .i_x2(w_pp_01_02),
    .i_x3(w_pp_02_01), .i_x4(w_pp_03_00),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_03_440), .ow_carry(w_c4to2_carry_03_440), .ow_cout(w_c4to2_cout_03_440)
);
wire w_c4to2_sum_04_441, w_c4to2_carry_04_441, w_c4to2_cout_04_441;
math_compressor_4to2 u_c4to2_04_441 (
    .i_x1(w_pp_04_00), .i_x2(w_c4to2_sum_04_360),
    .i_x3(w_c4to2_carry_03_440), .i_x4(w_c4to2_cout_03_440),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_04_441), .ow_carry(w_c4to2_carry_04_441), .ow_cout(w_c4to2_cout_04_441)
);
wire w_c4to2_sum_05_442, w_c4to2_carry_05_442, w_c4to2_cout_05_442;
math_compressor_4to2 u_c4to2_05_442 (
    .i_x1(w_c4to2_sum_05_361), .i_x2(w_c4to2_sum_05_362),
    .i_x3(w_c4to2_carry_04_441), .i_x4(w_c4to2_cout_04_441),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_05_442), .ow_carry(w_c4to2_carry_05_442), .ow_cout(w_c4to2_cout_05_442)
);
wire w_c4to2_sum_06_443, w_c4to2_carry_06_443, w_c4to2_cout_06_443;
math_compressor_4to2 u_c4to2_06_443 (
    .i_x1(w_c4to2_sum_06_363), .i_x2(w_c4to2_sum_06_364),
    .i_x3(w_c4to2_carry_05_442), .i_x4(w_c4to2_cout_05_442),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_06_443), .ow_carry(w_c4to2_carry_06_443), .ow_cout(w_c4to2_cout_06_443)
);
wire w_c4to2_sum_07_444, w_c4to2_carry_07_444, w_c4to2_cout_07_444;
math_compressor_4to2 u_c4to2_07_444 (
    .i_x1(w_c4to2_sum_07_365), .i_x2(w_c4to2_sum_07_366),
    .i_x3(w_c4to2_carry_06_443), .i_x4(w_c4to2_cout_06_443),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_07_444), .ow_carry(w_c4to2_carry_07_444), .ow_cout(w_c4to2_cout_07_444)
);
wire w_c4to2_sum_08_445, w_c4to2_carry_08_445, w_c4to2_cout_08_445;
math_compressor_4to2 u_c4to2_08_445 (
    .i_x1(w_c4to2_sum_08_367), .i_x2(w_c4to2_sum_08_368),
    .i_x3(w_c4to2_carry_07_444), .i_x4(w_c4to2_cout_07_444),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_08_445), .ow_carry(w_c4to2_carry_08_445), .ow_cout(w_c4to2_cout_08_445)
);
wire w_c4to2_sum_09_446, w_c4to2_carry_09_446, w_c4to2_cout_09_446;
math_compressor_4to2 u_c4to2_09_446 (
    .i_x1(w_c4to2_sum_09_369), .i_x2(w_c4to2_sum_09_370),
    .i_x3(w_c4to2_carry_08_445), .i_x4(w_c4to2_cout_08_445),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_09_446), .ow_carry(w_c4to2_carry_09_446), .ow_cout(w_c4to2_cout_09_446)
);
wire w_c4to2_sum_10_447, w_c4to2_carry_10_447, w_c4to2_cout_10_447;
math_compressor_4to2 u_c4to2_10_447 (
    .i_x1(w_c4to2_sum_10_371), .i_x2(w_c4to2_sum_10_372),
    .i_x3(w_c4to2_carry_09_446), .i_x4(w_c4to2_cout_09_446),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_10_447), .ow_carry(w_c4to2_carry_10_447), .ow_cout(w_c4to2_cout_10_447)
);
wire w_c4to2_sum_11_448, w_c4to2_carry_11_448, w_c4to2_cout_11_448;
math_compressor_4to2 u_c4to2_11_448 (
    .i_x1(w_c4to2_sum_11_373), .i_x2(w_c4to2_sum_11_374),
    .i_x3(w_c4to2_carry_10_447), .i_x4(w_c4to2_cout_10_447),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_11_448), .ow_carry(w_c4to2_carry_11_448), .ow_cout(w_c4to2_cout_11_448)
);
wire w_c4to2_sum_12_449, w_c4to2_carry_12_449, w_c4to2_cout_12_449;
math_compressor_4to2 u_c4to2_12_449 (
    .i_x1(w_c4to2_sum_12_375), .i_x2(w_c4to2_sum_12_376),
    .i_x3(w_c4to2_carry_11_448), .i_x4(w_c4to2_cout_11_448),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_12_449), .ow_carry(w_c4to2_carry_12_449), .ow_cout(w_c4to2_cout_12_449)
);
wire w_c4to2_sum_13_450, w_c4to2_carry_13_450, w_c4to2_cout_13_450;
math_compressor_4to2 u_c4to2_13_450 (
    .i_x1(w_c4to2_sum_13_377), .i_x2(w_c4to2_sum_13_378),
    .i_x3(w_c4to2_carry_12_449), .i_x4(w_c4to2_cout_12_449),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_13_450), .ow_carry(w_c4to2_carry_13_450), .ow_cout(w_c4to2_cout_13_450)
);
wire w_c4to2_sum_14_451, w_c4to2_carry_14_451, w_c4to2_cout_14_451;
math_compressor_4to2 u_c4to2_14_451 (
    .i_x1(w_c4to2_sum_14_379), .i_x2(w_c4to2_sum_14_380),
    .i_x3(w_c4to2_carry_13_450), .i_x4(w_c4to2_cout_13_450),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_14_451), .ow_carry(w_c4to2_carry_14_451), .ow_cout(w_c4to2_cout_14_451)
);
wire w_c4to2_sum_15_452, w_c4to2_carry_15_452, w_c4to2_cout_15_452;
math_compressor_4to2 u_c4to2_15_452 (
    .i_x1(w_c4to2_sum_15_381), .i_x2(w_c4to2_sum_15_382),
    .i_x3(w_c4to2_carry_14_451), .i_x4(w_c4to2_cout_14_451),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_15_452), .ow_carry(w_c4to2_carry_15_452), .ow_cout(w_c4to2_cout_15_452)
);
wire w_c4to2_sum_16_453, w_c4to2_carry_16_453, w_c4to2_cout_16_453;
math_compressor_4to2 u_c4to2_16_453 (
    .i_x1(w_c4to2_sum_16_383), .i_x2(w_c4to2_sum_16_384),
    .i_x3(w_c4to2_carry_15_452), .i_x4(w_c4to2_cout_15_452),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_16_453), .ow_carry(w_c4to2_carry_16_453), .ow_cout(w_c4to2_cout_16_453)
);
wire w_c4to2_sum_17_454, w_c4to2_carry_17_454, w_c4to2_cout_17_454;
math_compressor_4to2 u_c4to2_17_454 (
    .i_x1(w_c4to2_sum_17_385), .i_x2(w_c4to2_sum_17_386),
    .i_x3(w_c4to2_carry_16_453), .i_x4(w_c4to2_cout_16_453),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_17_454), .ow_carry(w_c4to2_carry_17_454), .ow_cout(w_c4to2_cout_17_454)
);
wire w_c4to2_sum_18_455, w_c4to2_carry_18_455, w_c4to2_cout_18_455;
math_compressor_4to2 u_c4to2_18_455 (
    .i_x1(w_c4to2_sum_18_387), .i_x2(w_c4to2_sum_18_388),
    .i_x3(w_c4to2_carry_17_454), .i_x4(w_c4to2_cout_17_454),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_18_455), .ow_carry(w_c4to2_carry_18_455), .ow_cout(w_c4to2_cout_18_455)
);
wire w_c4to2_sum_19_456, w_c4to2_carry_19_456, w_c4to2_cout_19_456;
math_compressor_4to2 u_c4to2_19_456 (
    .i_x1(w_c4to2_sum_19_389), .i_x2(w_c4to2_sum_19_390),
    .i_x3(w_c4to2_carry_18_455), .i_x4(w_c4to2_cout_18_455),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_19_456), .ow_carry(w_c4to2_carry_19_456), .ow_cout(w_c4to2_cout_19_456)
);
wire w_c4to2_sum_20_457, w_c4to2_carry_20_457, w_c4to2_cout_20_457;
math_compressor_4to2 u_c4to2_20_457 (
    .i_x1(w_c4to2_sum_20_391), .i_x2(w_c4to2_sum_20_392),
    .i_x3(w_c4to2_carry_19_456), .i_x4(w_c4to2_cout_19_456),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_20_457), .ow_carry(w_c4to2_carry_20_457), .ow_cout(w_c4to2_cout_20_457)
);
wire w_c4to2_sum_21_458, w_c4to2_carry_21_458, w_c4to2_cout_21_458;
math_compressor_4to2 u_c4to2_21_458 (
    .i_x1(w_c4to2_sum_21_393), .i_x2(w_c4to2_sum_21_394),
    .i_x3(w_c4to2_carry_20_457), .i_x4(w_c4to2_cout_20_457),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_21_458), .ow_carry(w_c4to2_carry_21_458), .ow_cout(w_c4to2_cout_21_458)
);
wire w_c4to2_sum_22_459, w_c4to2_carry_22_459, w_c4to2_cout_22_459;
math_compressor_4to2 u_c4to2_22_459 (
    .i_x1(w_c4to2_sum_22_395), .i_x2(w_c4to2_sum_22_396),
    .i_x3(w_c4to2_carry_21_458), .i_x4(w_c4to2_cout_21_458),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_22_459), .ow_carry(w_c4to2_carry_22_459), .ow_cout(w_c4to2_cout_22_459)
);
wire w_c4to2_sum_23_460, w_c4to2_carry_23_460, w_c4to2_cout_23_460;
math_compressor_4to2 u_c4to2_23_460 (
    .i_x1(w_c4to2_sum_23_397), .i_x2(w_c4to2_sum_23_398),
    .i_x3(w_c4to2_carry_22_459), .i_x4(w_c4to2_cout_22_459),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_23_460), .ow_carry(w_c4to2_carry_23_460), .ow_cout(w_c4to2_cout_23_460)
);
wire w_c4to2_sum_24_461, w_c4to2_carry_24_461, w_c4to2_cout_24_461;
math_compressor_4to2 u_c4to2_24_461 (
    .i_x1(w_c4to2_cout_23_398), .i_x2(w_c4to2_sum_24_399),
    .i_x3(w_c4to2_sum_24_400), .i_x4(w_c4to2_carry_23_460),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_24_461), .ow_carry(w_c4to2_carry_24_461), .ow_cout(w_c4to2_cout_24_461)
);
wire w_c4to2_sum_25_462, w_c4to2_carry_25_462, w_c4to2_cout_25_462;
math_compressor_4to2 u_c4to2_25_462 (
    .i_x1(w_c4to2_sum_25_401), .i_x2(w_c4to2_sum_25_402),
    .i_x3(w_c4to2_carry_24_461), .i_x4(w_c4to2_cout_24_461),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_25_462), .ow_carry(w_c4to2_carry_25_462), .ow_cout(w_c4to2_cout_25_462)
);
wire w_c4to2_sum_26_463, w_c4to2_carry_26_463, w_c4to2_cout_26_463;
math_compressor_4to2 u_c4to2_26_463 (
    .i_x1(w_c4to2_carry_25_402), .i_x2(w_c4to2_cout_25_402),
    .i_x3(w_c4to2_sum_26_403), .i_x4(w_c4to2_sum_26_404),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_26_463), .ow_carry(w_c4to2_carry_26_463), .ow_cout(w_c4to2_cout_26_463)
);
wire w_c4to2_sum_27_464, w_c4to2_carry_27_464, w_c4to2_cout_27_464;
math_compressor_4to2 u_c4to2_27_464 (
    .i_x1(w_c4to2_carry_26_404), .i_x2(w_c4to2_cout_26_404),
    .i_x3(w_c4to2_sum_27_405), .i_x4(w_c4to2_sum_27_406),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_464), .ow_carry(w_c4to2_carry_27_464), .ow_cout(w_c4to2_cout_27_464)
);
wire w_c4to2_sum_28_465, w_c4to2_carry_28_465, w_c4to2_cout_28_465;
math_compressor_4to2 u_c4to2_28_465 (
    .i_x1(w_c4to2_carry_27_406), .i_x2(w_c4to2_cout_27_406),
    .i_x3(w_c4to2_sum_28_407), .i_x4(w_c4to2_sum_28_408),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_465), .ow_carry(w_c4to2_carry_28_465), .ow_cout(w_c4to2_cout_28_465)
);
wire w_c4to2_sum_29_466, w_c4to2_carry_29_466, w_c4to2_cout_29_466;
math_compressor_4to2 u_c4to2_29_466 (
    .i_x1(w_c4to2_carry_28_408), .i_x2(w_c4to2_cout_28_408),
    .i_x3(w_c4to2_sum_29_409), .i_x4(w_c4to2_sum_29_410),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_466), .ow_carry(w_c4to2_carry_29_466), .ow_cout(w_c4to2_cout_29_466)
);
wire w_c4to2_sum_30_467, w_c4to2_carry_30_467, w_c4to2_cout_30_467;
math_compressor_4to2 u_c4to2_30_467 (
    .i_x1(w_c4to2_carry_29_410), .i_x2(w_c4to2_cout_29_410),
    .i_x3(w_c4to2_sum_30_411), .i_x4(w_c4to2_sum_30_412),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_467), .ow_carry(w_c4to2_carry_30_467), .ow_cout(w_c4to2_cout_30_467)
);
wire w_c4to2_sum_31_468, w_c4to2_carry_31_468, w_c4to2_cout_31_468;
math_compressor_4to2 u_c4to2_31_468 (
    .i_x1(w_c4to2_carry_30_412), .i_x2(w_c4to2_cout_30_412),
    .i_x3(w_c4to2_sum_31_413), .i_x4(w_c4to2_sum_31_414),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_468), .ow_carry(w_c4to2_carry_31_468), .ow_cout(w_c4to2_cout_31_468)
);
wire w_c4to2_sum_32_469, w_c4to2_carry_32_469, w_c4to2_cout_32_469;
math_compressor_4to2 u_c4to2_32_469 (
    .i_x1(w_c4to2_carry_31_414), .i_x2(w_c4to2_cout_31_414),
    .i_x3(w_c4to2_sum_32_415), .i_x4(w_c4to2_sum_32_416),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_469), .ow_carry(w_c4to2_carry_32_469), .ow_cout(w_c4to2_cout_32_469)
);
wire w_c4to2_sum_33_470, w_c4to2_carry_33_470, w_c4to2_cout_33_470;
math_compressor_4to2 u_c4to2_33_470 (
    .i_x1(w_c4to2_carry_32_416), .i_x2(w_c4to2_cout_32_416),
    .i_x3(w_c4to2_sum_33_417), .i_x4(w_c4to2_sum_33_418),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_470), .ow_carry(w_c4to2_carry_33_470), .ow_cout(w_c4to2_cout_33_470)
);
wire w_c4to2_sum_34_471, w_c4to2_carry_34_471, w_c4to2_cout_34_471;
math_compressor_4to2 u_c4to2_34_471 (
    .i_x1(w_c4to2_carry_33_418), .i_x2(w_c4to2_cout_33_418),
    .i_x3(w_c4to2_sum_34_419), .i_x4(w_c4to2_sum_34_420),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_471), .ow_carry(w_c4to2_carry_34_471), .ow_cout(w_c4to2_cout_34_471)
);
wire w_c4to2_sum_35_472, w_c4to2_carry_35_472, w_c4to2_cout_35_472;
math_compressor_4to2 u_c4to2_35_472 (
    .i_x1(w_c4to2_carry_34_420), .i_x2(w_c4to2_cout_34_420),
    .i_x3(w_c4to2_sum_35_421), .i_x4(w_c4to2_sum_35_422),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_472), .ow_carry(w_c4to2_carry_35_472), .ow_cout(w_c4to2_cout_35_472)
);
wire w_c4to2_sum_36_473, w_c4to2_carry_36_473, w_c4to2_cout_36_473;
math_compressor_4to2 u_c4to2_36_473 (
    .i_x1(w_c4to2_carry_35_422), .i_x2(w_c4to2_cout_35_422),
    .i_x3(w_c4to2_sum_36_423), .i_x4(w_c4to2_sum_36_424),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_473), .ow_carry(w_c4to2_carry_36_473), .ow_cout(w_c4to2_cout_36_473)
);
wire w_c4to2_sum_37_474, w_c4to2_carry_37_474, w_c4to2_cout_37_474;
math_compressor_4to2 u_c4to2_37_474 (
    .i_x1(w_c4to2_carry_36_424), .i_x2(w_c4to2_cout_36_424),
    .i_x3(w_c4to2_sum_37_425), .i_x4(w_c4to2_sum_37_426),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_474), .ow_carry(w_c4to2_carry_37_474), .ow_cout(w_c4to2_cout_37_474)
);
wire w_c4to2_sum_38_475, w_c4to2_carry_38_475, w_c4to2_cout_38_475;
math_compressor_4to2 u_c4to2_38_475 (
    .i_x1(w_c4to2_carry_37_426), .i_x2(w_c4to2_cout_37_426),
    .i_x3(w_c4to2_sum_38_427), .i_x4(w_c4to2_sum_38_428),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_475), .ow_carry(w_c4to2_carry_38_475), .ow_cout(w_c4to2_cout_38_475)
);
wire w_c4to2_sum_39_476, w_c4to2_carry_39_476, w_c4to2_cout_39_476;
math_compressor_4to2 u_c4to2_39_476 (
    .i_x1(w_c4to2_carry_38_428), .i_x2(w_c4to2_cout_38_428),
    .i_x3(w_c4to2_sum_39_429), .i_x4(w_c4to2_sum_39_430),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_476), .ow_carry(w_c4to2_carry_39_476), .ow_cout(w_c4to2_cout_39_476)
);
wire w_c4to2_sum_40_477, w_c4to2_carry_40_477, w_c4to2_cout_40_477;
math_compressor_4to2 u_c4to2_40_477 (
    .i_x1(w_c4to2_carry_39_430), .i_x2(w_c4to2_cout_39_430),
    .i_x3(w_c4to2_sum_40_431), .i_x4(w_c4to2_sum_40_432),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_477), .ow_carry(w_c4to2_carry_40_477), .ow_cout(w_c4to2_cout_40_477)
);
wire w_c4to2_sum_41_478, w_c4to2_carry_41_478, w_c4to2_cout_41_478;
math_compressor_4to2 u_c4to2_41_478 (
    .i_x1(w_c4to2_carry_40_432), .i_x2(w_c4to2_cout_40_432),
    .i_x3(w_c4to2_sum_41_433), .i_x4(w_c4to2_sum_41_434),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_478), .ow_carry(w_c4to2_carry_41_478), .ow_cout(w_c4to2_cout_41_478)
);
wire w_c4to2_sum_42_479, w_c4to2_carry_42_479, w_c4to2_cout_42_479;
math_compressor_4to2 u_c4to2_42_479 (
    .i_x1(w_c4to2_carry_41_434), .i_x2(w_c4to2_cout_41_434),
    .i_x3(w_c4to2_sum_42_435), .i_x4(w_c4to2_sum_42_436),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_42_479), .ow_carry(w_c4to2_carry_42_479), .ow_cout(w_c4to2_cout_42_479)
);
wire w_c4to2_sum_43_480, w_c4to2_carry_43_480, w_c4to2_cout_43_480;
math_compressor_4to2 u_c4to2_43_480 (
    .i_x1(w_c4to2_carry_42_436), .i_x2(w_c4to2_cout_42_436),
    .i_x3(w_c4to2_sum_43_437), .i_x4(w_c4to2_sum_43_438),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_43_480), .ow_carry(w_c4to2_carry_43_480), .ow_cout(w_c4to2_cout_43_480)
);
wire w_c4to2_sum_44_481, w_c4to2_carry_44_481, w_c4to2_cout_44_481;
math_compressor_4to2 u_c4to2_44_481 (
    .i_x1(w_c4to2_cout_43_437), .i_x2(w_c4to2_carry_43_438),
    .i_x3(w_c4to2_cout_43_438), .i_x4(w_c4to2_sum_44_439),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_44_481), .ow_carry(w_c4to2_carry_44_481), .ow_cout(w_c4to2_cout_44_481)
);
wire w_c4to2_sum_45_482, w_c4to2_carry_45_482, w_c4to2_cout_45_482;
math_compressor_4to2 u_c4to2_45_482 (
    .i_x1(w_pp_22_23), .i_x2(w_pp_23_22),
    .i_x3(w_c4to2_carry_44_439), .i_x4(w_c4to2_cout_44_439),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_45_482), .ow_carry(w_c4to2_carry_45_482), .ow_cout(w_c4to2_cout_45_482)
);

// Dadda Reduction Stage 7: height 3 -> 2

wire w_fa_sum_02_000, w_fa_carry_02_000;
math_adder_full u_fa_02_000 (
    .i_a(w_pp_00_02), .i_b(w_pp_01_01), .i_c(w_pp_02_00),
    .ow_sum(w_fa_sum_02_000), .ow_carry(w_fa_carry_02_000)
);
wire w_fa_sum_26_001, w_fa_carry_26_001;
math_adder_full u_fa_26_001 (
    .i_a(w_c4to2_carry_25_462), .i_b(w_c4to2_cout_25_462), .i_c(w_c4to2_sum_26_463),
    .ow_sum(w_fa_sum_26_001), .ow_carry(w_fa_carry_26_001)
);
wire w_c4to2_sum_27_483, w_c4to2_carry_27_483, w_c4to2_cout_27_483;
math_compressor_4to2 u_c4to2_27_483 (
    .i_x1(w_c4to2_carry_26_463), .i_x2(w_c4to2_cout_26_463),
    .i_x3(w_c4to2_sum_27_464), .i_x4(w_fa_carry_26_001),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_27_483), .ow_carry(w_c4to2_carry_27_483), .ow_cout(w_c4to2_cout_27_483)
);
wire w_c4to2_sum_28_484, w_c4to2_carry_28_484, w_c4to2_cout_28_484;
math_compressor_4to2 u_c4to2_28_484 (
    .i_x1(w_c4to2_carry_27_464), .i_x2(w_c4to2_cout_27_464),
    .i_x3(w_c4to2_sum_28_465), .i_x4(w_c4to2_carry_27_483),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_28_484), .ow_carry(w_c4to2_carry_28_484), .ow_cout(w_c4to2_cout_28_484)
);
wire w_c4to2_sum_29_485, w_c4to2_carry_29_485, w_c4to2_cout_29_485;
math_compressor_4to2 u_c4to2_29_485 (
    .i_x1(w_c4to2_carry_28_465), .i_x2(w_c4to2_cout_28_465),
    .i_x3(w_c4to2_sum_29_466), .i_x4(w_c4to2_carry_28_484),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_29_485), .ow_carry(w_c4to2_carry_29_485), .ow_cout(w_c4to2_cout_29_485)
);
wire w_c4to2_sum_30_486, w_c4to2_carry_30_486, w_c4to2_cout_30_486;
math_compressor_4to2 u_c4to2_30_486 (
    .i_x1(w_c4to2_carry_29_466), .i_x2(w_c4to2_cout_29_466),
    .i_x3(w_c4to2_sum_30_467), .i_x4(w_c4to2_carry_29_485),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_30_486), .ow_carry(w_c4to2_carry_30_486), .ow_cout(w_c4to2_cout_30_486)
);
wire w_c4to2_sum_31_487, w_c4to2_carry_31_487, w_c4to2_cout_31_487;
math_compressor_4to2 u_c4to2_31_487 (
    .i_x1(w_c4to2_carry_30_467), .i_x2(w_c4to2_cout_30_467),
    .i_x3(w_c4to2_sum_31_468), .i_x4(w_c4to2_carry_30_486),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_31_487), .ow_carry(w_c4to2_carry_31_487), .ow_cout(w_c4to2_cout_31_487)
);
wire w_c4to2_sum_32_488, w_c4to2_carry_32_488, w_c4to2_cout_32_488;
math_compressor_4to2 u_c4to2_32_488 (
    .i_x1(w_c4to2_carry_31_468), .i_x2(w_c4to2_cout_31_468),
    .i_x3(w_c4to2_sum_32_469), .i_x4(w_c4to2_carry_31_487),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_32_488), .ow_carry(w_c4to2_carry_32_488), .ow_cout(w_c4to2_cout_32_488)
);
wire w_c4to2_sum_33_489, w_c4to2_carry_33_489, w_c4to2_cout_33_489;
math_compressor_4to2 u_c4to2_33_489 (
    .i_x1(w_c4to2_carry_32_469), .i_x2(w_c4to2_cout_32_469),
    .i_x3(w_c4to2_sum_33_470), .i_x4(w_c4to2_carry_32_488),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_33_489), .ow_carry(w_c4to2_carry_33_489), .ow_cout(w_c4to2_cout_33_489)
);
wire w_c4to2_sum_34_490, w_c4to2_carry_34_490, w_c4to2_cout_34_490;
math_compressor_4to2 u_c4to2_34_490 (
    .i_x1(w_c4to2_carry_33_470), .i_x2(w_c4to2_cout_33_470),
    .i_x3(w_c4to2_sum_34_471), .i_x4(w_c4to2_carry_33_489),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_34_490), .ow_carry(w_c4to2_carry_34_490), .ow_cout(w_c4to2_cout_34_490)
);
wire w_c4to2_sum_35_491, w_c4to2_carry_35_491, w_c4to2_cout_35_491;
math_compressor_4to2 u_c4to2_35_491 (
    .i_x1(w_c4to2_carry_34_471), .i_x2(w_c4to2_cout_34_471),
    .i_x3(w_c4to2_sum_35_472), .i_x4(w_c4to2_carry_34_490),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_35_491), .ow_carry(w_c4to2_carry_35_491), .ow_cout(w_c4to2_cout_35_491)
);
wire w_c4to2_sum_36_492, w_c4to2_carry_36_492, w_c4to2_cout_36_492;
math_compressor_4to2 u_c4to2_36_492 (
    .i_x1(w_c4to2_carry_35_472), .i_x2(w_c4to2_cout_35_472),
    .i_x3(w_c4to2_sum_36_473), .i_x4(w_c4to2_carry_35_491),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_36_492), .ow_carry(w_c4to2_carry_36_492), .ow_cout(w_c4to2_cout_36_492)
);
wire w_c4to2_sum_37_493, w_c4to2_carry_37_493, w_c4to2_cout_37_493;
math_compressor_4to2 u_c4to2_37_493 (
    .i_x1(w_c4to2_carry_36_473), .i_x2(w_c4to2_cout_36_473),
    .i_x3(w_c4to2_sum_37_474), .i_x4(w_c4to2_carry_36_492),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_37_493), .ow_carry(w_c4to2_carry_37_493), .ow_cout(w_c4to2_cout_37_493)
);
wire w_c4to2_sum_38_494, w_c4to2_carry_38_494, w_c4to2_cout_38_494;
math_compressor_4to2 u_c4to2_38_494 (
    .i_x1(w_c4to2_carry_37_474), .i_x2(w_c4to2_cout_37_474),
    .i_x3(w_c4to2_sum_38_475), .i_x4(w_c4to2_carry_37_493),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_38_494), .ow_carry(w_c4to2_carry_38_494), .ow_cout(w_c4to2_cout_38_494)
);
wire w_c4to2_sum_39_495, w_c4to2_carry_39_495, w_c4to2_cout_39_495;
math_compressor_4to2 u_c4to2_39_495 (
    .i_x1(w_c4to2_carry_38_475), .i_x2(w_c4to2_cout_38_475),
    .i_x3(w_c4to2_sum_39_476), .i_x4(w_c4to2_carry_38_494),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_39_495), .ow_carry(w_c4to2_carry_39_495), .ow_cout(w_c4to2_cout_39_495)
);
wire w_c4to2_sum_40_496, w_c4to2_carry_40_496, w_c4to2_cout_40_496;
math_compressor_4to2 u_c4to2_40_496 (
    .i_x1(w_c4to2_carry_39_476), .i_x2(w_c4to2_cout_39_476),
    .i_x3(w_c4to2_sum_40_477), .i_x4(w_c4to2_carry_39_495),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_40_496), .ow_carry(w_c4to2_carry_40_496), .ow_cout(w_c4to2_cout_40_496)
);
wire w_c4to2_sum_41_497, w_c4to2_carry_41_497, w_c4to2_cout_41_497;
math_compressor_4to2 u_c4to2_41_497 (
    .i_x1(w_c4to2_carry_40_477), .i_x2(w_c4to2_cout_40_477),
    .i_x3(w_c4to2_sum_41_478), .i_x4(w_c4to2_carry_40_496),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_41_497), .ow_carry(w_c4to2_carry_41_497), .ow_cout(w_c4to2_cout_41_497)
);
wire w_c4to2_sum_42_498, w_c4to2_carry_42_498, w_c4to2_cout_42_498;
math_compressor_4to2 u_c4to2_42_498 (
    .i_x1(w_c4to2_carry_41_478), .i_x2(w_c4to2_cout_41_478),
    .i_x3(w_c4to2_sum_42_479), .i_x4(w_c4to2_carry_41_497),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_42_498), .ow_carry(w_c4to2_carry_42_498), .ow_cout(w_c4to2_cout_42_498)
);
wire w_c4to2_sum_43_499, w_c4to2_carry_43_499, w_c4to2_cout_43_499;
math_compressor_4to2 u_c4to2_43_499 (
    .i_x1(w_c4to2_carry_42_479), .i_x2(w_c4to2_cout_42_479),
    .i_x3(w_c4to2_sum_43_480), .i_x4(w_c4to2_carry_42_498),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_43_499), .ow_carry(w_c4to2_carry_43_499), .ow_cout(w_c4to2_cout_43_499)
);
wire w_c4to2_sum_44_500, w_c4to2_carry_44_500, w_c4to2_cout_44_500;
math_compressor_4to2 u_c4to2_44_500 (
    .i_x1(w_c4to2_carry_43_480), .i_x2(w_c4to2_cout_43_480),
    .i_x3(w_c4to2_sum_44_481), .i_x4(w_c4to2_carry_43_499),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_44_500), .ow_carry(w_c4to2_carry_44_500), .ow_cout(w_c4to2_cout_44_500)
);
wire w_c4to2_sum_45_501, w_c4to2_carry_45_501, w_c4to2_cout_45_501;
math_compressor_4to2 u_c4to2_45_501 (
    .i_x1(w_c4to2_carry_44_481), .i_x2(w_c4to2_cout_44_481),
    .i_x3(w_c4to2_sum_45_482), .i_x4(w_c4to2_carry_44_500),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_45_501), .ow_carry(w_c4to2_carry_45_501), .ow_cout(w_c4to2_cout_45_501)
);
wire w_c4to2_sum_46_502, w_c4to2_carry_46_502, w_c4to2_cout_46_502;
math_compressor_4to2 u_c4to2_46_502 (
    .i_x1(w_pp_23_23), .i_x2(w_c4to2_carry_45_482),
    .i_x3(w_c4to2_cout_45_482), .i_x4(w_c4to2_carry_45_501),
    .i_cin(1'b0),
    .ow_sum(w_c4to2_sum_46_502), .ow_carry(w_c4to2_carry_46_502), .ow_cout(w_c4to2_cout_46_502)
);

// Final CPA: Two operands from reduction tree
wire [2*N-1:0] w_cpa_a, w_cpa_b;
assign w_cpa_a[0] = w_pp_00_00;
assign w_cpa_b[0] = 1'b0;
assign w_cpa_a[1] = w_pp_00_01;
assign w_cpa_b[1] = w_pp_01_00;
assign w_cpa_a[2] = w_fa_sum_02_000;
assign w_cpa_b[2] = 1'b0;
assign w_cpa_a[3] = w_c4to2_sum_03_440;
assign w_cpa_b[3] = w_fa_carry_02_000;
assign w_cpa_a[4] = w_c4to2_sum_04_441;
assign w_cpa_b[4] = 1'b0;
assign w_cpa_a[5] = w_c4to2_sum_05_442;
assign w_cpa_b[5] = 1'b0;
assign w_cpa_a[6] = w_c4to2_sum_06_443;
assign w_cpa_b[6] = 1'b0;
assign w_cpa_a[7] = w_c4to2_sum_07_444;
assign w_cpa_b[7] = 1'b0;
assign w_cpa_a[8] = w_c4to2_sum_08_445;
assign w_cpa_b[8] = 1'b0;
assign w_cpa_a[9] = w_c4to2_sum_09_446;
assign w_cpa_b[9] = 1'b0;
assign w_cpa_a[10] = w_c4to2_sum_10_447;
assign w_cpa_b[10] = 1'b0;
assign w_cpa_a[11] = w_c4to2_sum_11_448;
assign w_cpa_b[11] = 1'b0;
assign w_cpa_a[12] = w_c4to2_sum_12_449;
assign w_cpa_b[12] = 1'b0;
assign w_cpa_a[13] = w_c4to2_sum_13_450;
assign w_cpa_b[13] = 1'b0;
assign w_cpa_a[14] = w_c4to2_sum_14_451;
assign w_cpa_b[14] = 1'b0;
assign w_cpa_a[15] = w_c4to2_sum_15_452;
assign w_cpa_b[15] = 1'b0;
assign w_cpa_a[16] = w_c4to2_sum_16_453;
assign w_cpa_b[16] = 1'b0;
assign w_cpa_a[17] = w_c4to2_sum_17_454;
assign w_cpa_b[17] = 1'b0;
assign w_cpa_a[18] = w_c4to2_sum_18_455;
assign w_cpa_b[18] = 1'b0;
assign w_cpa_a[19] = w_c4to2_sum_19_456;
assign w_cpa_b[19] = 1'b0;
assign w_cpa_a[20] = w_c4to2_sum_20_457;
assign w_cpa_b[20] = 1'b0;
assign w_cpa_a[21] = w_c4to2_sum_21_458;
assign w_cpa_b[21] = 1'b0;
assign w_cpa_a[22] = w_c4to2_sum_22_459;
assign w_cpa_b[22] = 1'b0;
assign w_cpa_a[23] = w_c4to2_sum_23_460;
assign w_cpa_b[23] = 1'b0;
assign w_cpa_a[24] = w_c4to2_cout_23_460;
assign w_cpa_b[24] = w_c4to2_sum_24_461;
assign w_cpa_a[25] = w_c4to2_sum_25_462;
assign w_cpa_b[25] = 1'b0;
assign w_cpa_a[26] = w_fa_sum_26_001;
assign w_cpa_b[26] = 1'b0;
assign w_cpa_a[27] = w_c4to2_sum_27_483;
assign w_cpa_b[27] = 1'b0;
assign w_cpa_a[28] = w_c4to2_cout_27_483;
assign w_cpa_b[28] = w_c4to2_sum_28_484;
assign w_cpa_a[29] = w_c4to2_cout_28_484;
assign w_cpa_b[29] = w_c4to2_sum_29_485;
assign w_cpa_a[30] = w_c4to2_cout_29_485;
assign w_cpa_b[30] = w_c4to2_sum_30_486;
assign w_cpa_a[31] = w_c4to2_cout_30_486;
assign w_cpa_b[31] = w_c4to2_sum_31_487;
assign w_cpa_a[32] = w_c4to2_cout_31_487;
assign w_cpa_b[32] = w_c4to2_sum_32_488;
assign w_cpa_a[33] = w_c4to2_cout_32_488;
assign w_cpa_b[33] = w_c4to2_sum_33_489;
assign w_cpa_a[34] = w_c4to2_cout_33_489;
assign w_cpa_b[34] = w_c4to2_sum_34_490;
assign w_cpa_a[35] = w_c4to2_cout_34_490;
assign w_cpa_b[35] = w_c4to2_sum_35_491;
assign w_cpa_a[36] = w_c4to2_cout_35_491;
assign w_cpa_b[36] = w_c4to2_sum_36_492;
assign w_cpa_a[37] = w_c4to2_cout_36_492;
assign w_cpa_b[37] = w_c4to2_sum_37_493;
assign w_cpa_a[38] = w_c4to2_cout_37_493;
assign w_cpa_b[38] = w_c4to2_sum_38_494;
assign w_cpa_a[39] = w_c4to2_cout_38_494;
assign w_cpa_b[39] = w_c4to2_sum_39_495;
assign w_cpa_a[40] = w_c4to2_cout_39_495;
assign w_cpa_b[40] = w_c4to2_sum_40_496;
assign w_cpa_a[41] = w_c4to2_cout_40_496;
assign w_cpa_b[41] = w_c4to2_sum_41_497;
assign w_cpa_a[42] = w_c4to2_cout_41_497;
assign w_cpa_b[42] = w_c4to2_sum_42_498;
assign w_cpa_a[43] = w_c4to2_cout_42_498;
assign w_cpa_b[43] = w_c4to2_sum_43_499;
assign w_cpa_a[44] = w_c4to2_cout_43_499;
assign w_cpa_b[44] = w_c4to2_sum_44_500;
assign w_cpa_a[45] = w_c4to2_cout_44_500;
assign w_cpa_b[45] = w_c4to2_sum_45_501;
assign w_cpa_a[46] = w_c4to2_cout_45_501;
assign w_cpa_b[46] = w_c4to2_sum_46_502;
assign w_cpa_a[47] = w_c4to2_carry_46_502;
assign w_cpa_b[47] = w_c4to2_cout_46_502;

// Han-Carlson prefix adder for final CPA
wire w_cpa_cout;  // Unused for unsigned multiply
math_adder_han_carlson_048 u_final_cpa (
    .i_a(w_cpa_a),
    .i_b(w_cpa_b),
    .i_cin(1'b0),
    .ow_sum(ow_product),
    .ow_cout(w_cpa_cout)
);

endmodule
