`timescale 1ns / 1ps

module math_multiplier_wallace_tree_csa_8 (
    input  [7:0] i_multiplier,
    input  [7:0] i_multiplicand,
    output [15:0] ow_product
);

// Partial products generation
wire w_pp_0_0 = i_multiplier[0] & i_multiplicand[0];
wire w_pp_0_1 = i_multiplier[0] & i_multiplicand[1];
wire w_pp_0_2 = i_multiplier[0] & i_multiplicand[2];
wire w_pp_0_3 = i_multiplier[0] & i_multiplicand[3];
wire w_pp_0_4 = i_multiplier[0] & i_multiplicand[4];
wire w_pp_0_5 = i_multiplier[0] & i_multiplicand[5];
wire w_pp_0_6 = i_multiplier[0] & i_multiplicand[6];
wire w_pp_0_7 = i_multiplier[0] & i_multiplicand[7];
wire w_pp_1_0 = i_multiplier[1] & i_multiplicand[0];
wire w_pp_1_1 = i_multiplier[1] & i_multiplicand[1];
wire w_pp_1_2 = i_multiplier[1] & i_multiplicand[2];
wire w_pp_1_3 = i_multiplier[1] & i_multiplicand[3];
wire w_pp_1_4 = i_multiplier[1] & i_multiplicand[4];
wire w_pp_1_5 = i_multiplier[1] & i_multiplicand[5];
wire w_pp_1_6 = i_multiplier[1] & i_multiplicand[6];
wire w_pp_1_7 = i_multiplier[1] & i_multiplicand[7];
wire w_pp_2_0 = i_multiplier[2] & i_multiplicand[0];
wire w_pp_2_1 = i_multiplier[2] & i_multiplicand[1];
wire w_pp_2_2 = i_multiplier[2] & i_multiplicand[2];
wire w_pp_2_3 = i_multiplier[2] & i_multiplicand[3];
wire w_pp_2_4 = i_multiplier[2] & i_multiplicand[4];
wire w_pp_2_5 = i_multiplier[2] & i_multiplicand[5];
wire w_pp_2_6 = i_multiplier[2] & i_multiplicand[6];
wire w_pp_2_7 = i_multiplier[2] & i_multiplicand[7];
wire w_pp_3_0 = i_multiplier[3] & i_multiplicand[0];
wire w_pp_3_1 = i_multiplier[3] & i_multiplicand[1];
wire w_pp_3_2 = i_multiplier[3] & i_multiplicand[2];
wire w_pp_3_3 = i_multiplier[3] & i_multiplicand[3];
wire w_pp_3_4 = i_multiplier[3] & i_multiplicand[4];
wire w_pp_3_5 = i_multiplier[3] & i_multiplicand[5];
wire w_pp_3_6 = i_multiplier[3] & i_multiplicand[6];
wire w_pp_3_7 = i_multiplier[3] & i_multiplicand[7];
wire w_pp_4_0 = i_multiplier[4] & i_multiplicand[0];
wire w_pp_4_1 = i_multiplier[4] & i_multiplicand[1];
wire w_pp_4_2 = i_multiplier[4] & i_multiplicand[2];
wire w_pp_4_3 = i_multiplier[4] & i_multiplicand[3];
wire w_pp_4_4 = i_multiplier[4] & i_multiplicand[4];
wire w_pp_4_5 = i_multiplier[4] & i_multiplicand[5];
wire w_pp_4_6 = i_multiplier[4] & i_multiplicand[6];
wire w_pp_4_7 = i_multiplier[4] & i_multiplicand[7];
wire w_pp_5_0 = i_multiplier[5] & i_multiplicand[0];
wire w_pp_5_1 = i_multiplier[5] & i_multiplicand[1];
wire w_pp_5_2 = i_multiplier[5] & i_multiplicand[2];
wire w_pp_5_3 = i_multiplier[5] & i_multiplicand[3];
wire w_pp_5_4 = i_multiplier[5] & i_multiplicand[4];
wire w_pp_5_5 = i_multiplier[5] & i_multiplicand[5];
wire w_pp_5_6 = i_multiplier[5] & i_multiplicand[6];
wire w_pp_5_7 = i_multiplier[5] & i_multiplicand[7];
wire w_pp_6_0 = i_multiplier[6] & i_multiplicand[0];
wire w_pp_6_1 = i_multiplier[6] & i_multiplicand[1];
wire w_pp_6_2 = i_multiplier[6] & i_multiplicand[2];
wire w_pp_6_3 = i_multiplier[6] & i_multiplicand[3];
wire w_pp_6_4 = i_multiplier[6] & i_multiplicand[4];
wire w_pp_6_5 = i_multiplier[6] & i_multiplicand[5];
wire w_pp_6_6 = i_multiplier[6] & i_multiplicand[6];
wire w_pp_6_7 = i_multiplier[6] & i_multiplicand[7];
wire w_pp_7_0 = i_multiplier[7] & i_multiplicand[0];
wire w_pp_7_1 = i_multiplier[7] & i_multiplicand[1];
wire w_pp_7_2 = i_multiplier[7] & i_multiplicand[2];
wire w_pp_7_3 = i_multiplier[7] & i_multiplicand[3];
wire w_pp_7_4 = i_multiplier[7] & i_multiplicand[4];
wire w_pp_7_5 = i_multiplier[7] & i_multiplicand[5];
wire w_pp_7_6 = i_multiplier[7] & i_multiplicand[6];
wire w_pp_7_7 = i_multiplier[7] & i_multiplicand[7];

// Partial products reduction using Wallace tree
wire w_sum_1_2, w_carry_1_2;
math_adder_half HA_1_2(.i_a(w_pp_0_1), .i_b(w_pp_1_0), .ow_sum(w_sum_1_2), .ow_c(w_carry_1_2));
wire w_sum_2_4, w_carry_2_4;
math_adder_carry_save CSA_2_4(.i_a(w_pp_0_2), .i_b(w_pp_1_1), .i_c(w_pp_2_0), .ow_sum(w_sum_2_4), .ow_c(w_carry_2_4));
wire w_sum_2_2, w_carry_2_2;
math_adder_half HA_2_2(.i_a(w_carry_1_2), .i_b(w_sum_2_4), .ow_sum(w_sum_2_2), .ow_c(w_carry_2_2));
wire w_sum_3_6, w_carry_3_6;
math_adder_carry_save CSA_3_6(.i_a(w_pp_0_3), .i_b(w_pp_1_2), .i_c(w_pp_2_1), .ow_sum(w_sum_3_6), .ow_c(w_carry_3_6));
wire w_sum_3_4, w_carry_3_4;
math_adder_carry_save CSA_3_4(.i_a(w_pp_3_0), .i_b(w_carry_2_4), .i_c(w_carry_2_2), .ow_sum(w_sum_3_4), .ow_c(w_carry_3_4));
wire w_sum_3_2, w_carry_3_2;
math_adder_half HA_3_2(.i_a(w_sum_3_6), .i_b(w_sum_3_4), .ow_sum(w_sum_3_2), .ow_c(w_carry_3_2));
wire w_sum_4_8, w_carry_4_8;
math_adder_carry_save CSA_4_8(.i_a(w_pp_0_4), .i_b(w_pp_1_3), .i_c(w_pp_2_2), .ow_sum(w_sum_4_8), .ow_c(w_carry_4_8));
wire w_sum_4_6, w_carry_4_6;
math_adder_carry_save CSA_4_6(.i_a(w_pp_3_1), .i_b(w_pp_4_0), .i_c(w_carry_3_6), .ow_sum(w_sum_4_6), .ow_c(w_carry_4_6));
wire w_sum_4_4, w_carry_4_4;
math_adder_carry_save CSA_4_4(.i_a(w_carry_3_4), .i_b(w_carry_3_2), .i_c(w_sum_4_8), .ow_sum(w_sum_4_4), .ow_c(w_carry_4_4));
wire w_sum_4_2, w_carry_4_2;
math_adder_half HA_4_2(.i_a(w_sum_4_6), .i_b(w_sum_4_4), .ow_sum(w_sum_4_2), .ow_c(w_carry_4_2));
wire w_sum_5_10, w_carry_5_10;
math_adder_carry_save CSA_5_10(.i_a(w_pp_0_5), .i_b(w_pp_1_4), .i_c(w_pp_2_3), .ow_sum(w_sum_5_10), .ow_c(w_carry_5_10));
wire w_sum_5_8, w_carry_5_8;
math_adder_carry_save CSA_5_8(.i_a(w_pp_3_2), .i_b(w_pp_4_1), .i_c(w_pp_5_0), .ow_sum(w_sum_5_8), .ow_c(w_carry_5_8));
wire w_sum_5_6, w_carry_5_6;
math_adder_carry_save CSA_5_6(.i_a(w_carry_4_8), .i_b(w_carry_4_6), .i_c(w_carry_4_4), .ow_sum(w_sum_5_6), .ow_c(w_carry_5_6));
wire w_sum_5_4, w_carry_5_4;
math_adder_carry_save CSA_5_4(.i_a(w_carry_4_2), .i_b(w_sum_5_10), .i_c(w_sum_5_8), .ow_sum(w_sum_5_4), .ow_c(w_carry_5_4));
wire w_sum_5_2, w_carry_5_2;
math_adder_half HA_5_2(.i_a(w_sum_5_6), .i_b(w_sum_5_4), .ow_sum(w_sum_5_2), .ow_c(w_carry_5_2));
wire w_sum_6_12, w_carry_6_12;
math_adder_carry_save CSA_6_12(.i_a(w_pp_0_6), .i_b(w_pp_1_5), .i_c(w_pp_2_4), .ow_sum(w_sum_6_12), .ow_c(w_carry_6_12));
wire w_sum_6_10, w_carry_6_10;
math_adder_carry_save CSA_6_10(.i_a(w_pp_3_3), .i_b(w_pp_4_2), .i_c(w_pp_5_1), .ow_sum(w_sum_6_10), .ow_c(w_carry_6_10));
wire w_sum_6_8, w_carry_6_8;
math_adder_carry_save CSA_6_8(.i_a(w_pp_6_0), .i_b(w_carry_5_10), .i_c(w_carry_5_8), .ow_sum(w_sum_6_8), .ow_c(w_carry_6_8));
wire w_sum_6_6, w_carry_6_6;
math_adder_carry_save CSA_6_6(.i_a(w_carry_5_6), .i_b(w_carry_5_4), .i_c(w_carry_5_2), .ow_sum(w_sum_6_6), .ow_c(w_carry_6_6));
wire w_sum_6_4, w_carry_6_4;
math_adder_carry_save CSA_6_4(.i_a(w_sum_6_12), .i_b(w_sum_6_10), .i_c(w_sum_6_8), .ow_sum(w_sum_6_4), .ow_c(w_carry_6_4));
wire w_sum_6_2, w_carry_6_2;
math_adder_half HA_6_2(.i_a(w_sum_6_6), .i_b(w_sum_6_4), .ow_sum(w_sum_6_2), .ow_c(w_carry_6_2));
wire w_sum_7_14, w_carry_7_14;
math_adder_carry_save CSA_7_14(.i_a(w_pp_0_7), .i_b(w_pp_1_6), .i_c(w_pp_2_5), .ow_sum(w_sum_7_14), .ow_c(w_carry_7_14));
wire w_sum_7_12, w_carry_7_12;
math_adder_carry_save CSA_7_12(.i_a(w_pp_3_4), .i_b(w_pp_4_3), .i_c(w_pp_5_2), .ow_sum(w_sum_7_12), .ow_c(w_carry_7_12));
wire w_sum_7_10, w_carry_7_10;
math_adder_carry_save CSA_7_10(.i_a(w_pp_6_1), .i_b(w_pp_7_0), .i_c(w_carry_6_12), .ow_sum(w_sum_7_10), .ow_c(w_carry_7_10));
wire w_sum_7_8, w_carry_7_8;
math_adder_carry_save CSA_7_8(.i_a(w_carry_6_10), .i_b(w_carry_6_8), .i_c(w_carry_6_6), .ow_sum(w_sum_7_8), .ow_c(w_carry_7_8));
wire w_sum_7_6, w_carry_7_6;
math_adder_carry_save CSA_7_6(.i_a(w_carry_6_4), .i_b(w_carry_6_2), .i_c(w_sum_7_14), .ow_sum(w_sum_7_6), .ow_c(w_carry_7_6));
wire w_sum_7_4, w_carry_7_4;
math_adder_carry_save CSA_7_4(.i_a(w_sum_7_12), .i_b(w_sum_7_10), .i_c(w_sum_7_8), .ow_sum(w_sum_7_4), .ow_c(w_carry_7_4));
wire w_sum_7_2, w_carry_7_2;
math_adder_half HA_7_2(.i_a(w_sum_7_6), .i_b(w_sum_7_4), .ow_sum(w_sum_7_2), .ow_c(w_carry_7_2));
wire w_sum_8_14, w_carry_8_14;
math_adder_carry_save CSA_8_14(.i_a(w_pp_1_7), .i_b(w_pp_2_6), .i_c(w_pp_3_5), .ow_sum(w_sum_8_14), .ow_c(w_carry_8_14));
wire w_sum_8_12, w_carry_8_12;
math_adder_carry_save CSA_8_12(.i_a(w_pp_4_4), .i_b(w_pp_5_3), .i_c(w_pp_6_2), .ow_sum(w_sum_8_12), .ow_c(w_carry_8_12));
wire w_sum_8_10, w_carry_8_10;
math_adder_carry_save CSA_8_10(.i_a(w_pp_7_1), .i_b(w_carry_7_14), .i_c(w_carry_7_12), .ow_sum(w_sum_8_10), .ow_c(w_carry_8_10));
wire w_sum_8_8, w_carry_8_8;
math_adder_carry_save CSA_8_8(.i_a(w_carry_7_10), .i_b(w_carry_7_8), .i_c(w_carry_7_6), .ow_sum(w_sum_8_8), .ow_c(w_carry_8_8));
wire w_sum_8_6, w_carry_8_6;
math_adder_carry_save CSA_8_6(.i_a(w_carry_7_4), .i_b(w_carry_7_2), .i_c(w_sum_8_14), .ow_sum(w_sum_8_6), .ow_c(w_carry_8_6));
wire w_sum_8_4, w_carry_8_4;
math_adder_carry_save CSA_8_4(.i_a(w_sum_8_12), .i_b(w_sum_8_10), .i_c(w_sum_8_8), .ow_sum(w_sum_8_4), .ow_c(w_carry_8_4));
wire w_sum_8_2, w_carry_8_2;
math_adder_half HA_8_2(.i_a(w_sum_8_6), .i_b(w_sum_8_4), .ow_sum(w_sum_8_2), .ow_c(w_carry_8_2));
wire w_sum_9_13, w_carry_9_13;
math_adder_carry_save CSA_9_13(.i_a(w_pp_2_7), .i_b(w_pp_3_6), .i_c(w_pp_4_5), .ow_sum(w_sum_9_13), .ow_c(w_carry_9_13));
wire w_sum_9_11, w_carry_9_11;
math_adder_carry_save CSA_9_11(.i_a(w_pp_5_4), .i_b(w_pp_6_3), .i_c(w_pp_7_2), .ow_sum(w_sum_9_11), .ow_c(w_carry_9_11));
wire w_sum_9_9, w_carry_9_9;
math_adder_carry_save CSA_9_9(.i_a(w_carry_8_14), .i_b(w_carry_8_12), .i_c(w_carry_8_10), .ow_sum(w_sum_9_9), .ow_c(w_carry_9_9));
wire w_sum_9_7, w_carry_9_7;
math_adder_carry_save CSA_9_7(.i_a(w_carry_8_8), .i_b(w_carry_8_6), .i_c(w_carry_8_4), .ow_sum(w_sum_9_7), .ow_c(w_carry_9_7));
wire w_sum_9_5, w_carry_9_5;
math_adder_carry_save CSA_9_5(.i_a(w_carry_8_2), .i_b(w_sum_9_13), .i_c(w_sum_9_11), .ow_sum(w_sum_9_5), .ow_c(w_carry_9_5));
wire w_sum_9_3, w_carry_9_3;
math_adder_carry_save CSA_9_3(.i_a(w_sum_9_9), .i_b(w_sum_9_7), .i_c(w_sum_9_5), .ow_sum(w_sum_9_3), .ow_c(w_carry_9_3));
wire w_sum_10_11, w_carry_10_11;
math_adder_carry_save CSA_10_11(.i_a(w_pp_3_7), .i_b(w_pp_4_6), .i_c(w_pp_5_5), .ow_sum(w_sum_10_11), .ow_c(w_carry_10_11));
wire w_sum_10_9, w_carry_10_9;
math_adder_carry_save CSA_10_9(.i_a(w_pp_6_4), .i_b(w_pp_7_3), .i_c(w_carry_9_13), .ow_sum(w_sum_10_9), .ow_c(w_carry_10_9));
wire w_sum_10_7, w_carry_10_7;
math_adder_carry_save CSA_10_7(.i_a(w_carry_9_11), .i_b(w_carry_9_9), .i_c(w_carry_9_7), .ow_sum(w_sum_10_7), .ow_c(w_carry_10_7));
wire w_sum_10_5, w_carry_10_5;
math_adder_carry_save CSA_10_5(.i_a(w_carry_9_5), .i_b(w_carry_9_3), .i_c(w_sum_10_11), .ow_sum(w_sum_10_5), .ow_c(w_carry_10_5));
wire w_sum_10_3, w_carry_10_3;
math_adder_carry_save CSA_10_3(.i_a(w_sum_10_9), .i_b(w_sum_10_7), .i_c(w_sum_10_5), .ow_sum(w_sum_10_3), .ow_c(w_carry_10_3));
wire w_sum_11_9, w_carry_11_9;
math_adder_carry_save CSA_11_9(.i_a(w_pp_4_7), .i_b(w_pp_5_6), .i_c(w_pp_6_5), .ow_sum(w_sum_11_9), .ow_c(w_carry_11_9));
wire w_sum_11_7, w_carry_11_7;
math_adder_carry_save CSA_11_7(.i_a(w_pp_7_4), .i_b(w_carry_10_11), .i_c(w_carry_10_9), .ow_sum(w_sum_11_7), .ow_c(w_carry_11_7));
wire w_sum_11_5, w_carry_11_5;
math_adder_carry_save CSA_11_5(.i_a(w_carry_10_7), .i_b(w_carry_10_5), .i_c(w_carry_10_3), .ow_sum(w_sum_11_5), .ow_c(w_carry_11_5));
wire w_sum_11_3, w_carry_11_3;
math_adder_carry_save CSA_11_3(.i_a(w_sum_11_9), .i_b(w_sum_11_7), .i_c(w_sum_11_5), .ow_sum(w_sum_11_3), .ow_c(w_carry_11_3));
wire w_sum_12_7, w_carry_12_7;
math_adder_carry_save CSA_12_7(.i_a(w_pp_5_7), .i_b(w_pp_6_6), .i_c(w_pp_7_5), .ow_sum(w_sum_12_7), .ow_c(w_carry_12_7));
wire w_sum_12_5, w_carry_12_5;
math_adder_carry_save CSA_12_5(.i_a(w_carry_11_9), .i_b(w_carry_11_7), .i_c(w_carry_11_5), .ow_sum(w_sum_12_5), .ow_c(w_carry_12_5));
wire w_sum_12_3, w_carry_12_3;
math_adder_carry_save CSA_12_3(.i_a(w_carry_11_3), .i_b(w_sum_12_7), .i_c(w_sum_12_5), .ow_sum(w_sum_12_3), .ow_c(w_carry_12_3));
wire w_sum_13_5, w_carry_13_5;
math_adder_carry_save CSA_13_5(.i_a(w_pp_6_7), .i_b(w_pp_7_6), .i_c(w_carry_12_7), .ow_sum(w_sum_13_5), .ow_c(w_carry_13_5));
wire w_sum_13_3, w_carry_13_3;
math_adder_carry_save CSA_13_3(.i_a(w_carry_12_5), .i_b(w_carry_12_3), .i_c(w_sum_13_5), .ow_sum(w_sum_13_3), .ow_c(w_carry_13_3));
wire w_sum_14_3, w_carry_14_3;
math_adder_carry_save CSA_14_3(.i_a(w_pp_7_7), .i_b(w_carry_13_5), .i_c(w_carry_13_3), .ow_sum(w_sum_14_3), .ow_c(w_carry_14_3));

// Final product assignment
assign ow_product[0] = w_pp_0_0;
assign ow_product[1] = w_sum_1_2;
assign ow_product[2] = w_sum_2_2;
assign ow_product[3] = w_sum_3_2;
assign ow_product[4] = w_sum_4_2;
assign ow_product[5] = w_sum_5_2;
assign ow_product[6] = w_sum_6_2;
assign ow_product[7] = w_sum_7_2;
assign ow_product[8] = w_sum_8_2;
assign ow_product[9] = w_sum_9_3;
assign ow_product[10] = w_sum_10_3;
assign ow_product[11] = w_sum_11_3;
assign ow_product[12] = w_sum_12_3;
assign ow_product[13] = w_sum_13_3;
assign ow_product[14] = w_sum_14_3;
assign ow_product[15] = w_carry_14_3;


    // Debug purposes
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_wallace_tree_csa_8);
    end
                
endmodule : math_multiplier_wallace_tree_csa_8
