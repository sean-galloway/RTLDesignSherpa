// SPDX-License-Identifier: MIT
// SPDX-FileCopyrightText: 2024-2025 sean galloway
//
// RTL Design Sherpa - Industry-Standard RTL Design and Verification
// https://github.com/sean-galloway/RTLDesignSherpa
//
// Module: delta_axis_flat_3x8
// Purpose: AXI-Stream 3×8 Flat Crossbar Switch
//
// Documentation: projects/components/delta/PRD.md
// Subsystem: delta
//
// Author: sean galloway
// Created: 2025-10-18

`timescale 1ns / 1ps

module delta_axis_flat_3x8 #(parameter int  DATA_WIDTH = 64,
parameter int  DEST_WIDTH = 3,
parameter int  ID_WIDTH = 2,
parameter int  USER_WIDTH = 1,
parameter int  NUM_MASTERS = 3,
parameter int  NUM_SLAVES = 8 )(
    input  logic                  aclk,
    input  logic                  aresetn,
    input  logic [DATA_WIDTH-1:0] s_axis_tdata  [NUM_MASTERS],
    input  logic                  s_axis_tvalid [NUM_MASTERS],
    output logic                  s_axis_tready [NUM_MASTERS],
    input  logic                  s_axis_tlast  [NUM_MASTERS],
    input  logic [DEST_WIDTH-1:0] s_axis_tdest  [NUM_MASTERS],
    input  logic [ID_WIDTH-1:0]   s_axis_tid    [NUM_MASTERS],
    input  logic [USER_WIDTH-1:0] s_axis_tuser  [NUM_MASTERS],
    output logic [DATA_WIDTH-1:0] m_axis_tdata  [NUM_SLAVES],
    output logic                  m_axis_tvalid [NUM_SLAVES],
    input  logic                  m_axis_tready [NUM_SLAVES],
    output logic                  m_axis_tlast  [NUM_SLAVES],
    output logic [DEST_WIDTH-1:0] m_axis_tdest  [NUM_SLAVES],
    output logic [ID_WIDTH-1:0]   m_axis_tid    [NUM_SLAVES],
    output logic [USER_WIDTH-1:0] m_axis_tuser  [NUM_SLAVES]
);

// ==============================================================================
// Module: delta_axis_flat_3x8
// Project: Delta - AXI-Stream Crossbar Generator
// ==============================================================================
// Description: AXI-Stream 3×8 Flat Crossbar Switch
// 
// Delta: Where data flows split and merge like river deltas
// 
// Generated by: delta_generator_v2.py (framework version)
// Configuration:
//   - Topology: flat
//   - Masters: 3
//   - Slaves: 8
//   - Data Width: 64 bits
//   - TDEST Width: 3 bits
//   - TID Width: 2 bits
//   - Arbiter: round_robin
// 
// Features:
//   - Per-slave round-robin arbitration
//   - Packet atomicity (locked grant until TLAST)
//   - Registered outputs for timing closure
//   - Full AXI-Stream compliance
// 
// ==============================================================================

// ==========================================================================
// Request Generation - Decode TDEST to slave select
// ==========================================================================
// AXIS Advantage: Direct TDEST decode (simpler than APB address ranges)
// 
// Each master's TDEST field directly identifies target slave
// No address range checking needed (unlike APB crossbar)
// ==========================================================================

logic [NUM_MASTERS-1:0] request_matrix [NUM_SLAVES];

always_comb begin
    // Initialize all requests to zero
    for (int s = 0; s < NUM_SLAVES; s++) begin
        request_matrix[s] = '0;
    end

    // Generate requests based on TDEST
    for (int m = 0; m < NUM_MASTERS; m++) begin
        if (s_axis_tvalid[m] && (s_axis_tdest[m] < NUM_SLAVES[$clog2(NUM_SLAVES+1)-1:0])) begin
            // Direct decode: TDEST is slave index
            request_matrix[s_axis_tdest[m]][m] = 1'b1;
        end
    end
end

// ==========================================================================
// Per-Slave Round-Robin Arbiters with Packet Atomicity
// ==========================================================================
// Similar to APB crossbar, but with PACKET ATOMICITY:
// - APB: Re-arbitrate every cycle
// - AXIS: Lock grant until TLAST (prevent packet interleaving)
// 
// Round-robin ensures fair bandwidth allocation
// Packet atomicity ensures correct streaming behavior
// ==========================================================================

logic [NUM_MASTERS-1:0] grant_matrix [NUM_SLAVES];
logic [$clog2(NUM_MASTERS)-1:0] last_grant [NUM_SLAVES];
logic packet_active [NUM_SLAVES];  // NEW vs APB: Track packet in progress

// Arbitration logic for each slave
generate
    for (genvar s = 0; s < NUM_SLAVES; s++) begin : gen_arbiter
        always_ff @(posedge aclk or negedge aresetn) begin
            if (!aresetn) begin
                grant_matrix[s] <= '0;
                last_grant[s] <= '0;
                packet_active[s] <= 1'b0;
            end else begin
                if (packet_active[s]) begin
                    // Hold grant until TLAST (packet atomicity)
                    if (m_axis_tvalid[s] && m_axis_tready[s] && m_axis_tlast[s]) begin
                        packet_active[s] <= 1'b0;
                        grant_matrix[s] <= '0;
                    end
                end else if (|request_matrix[s]) begin
                    // Round-robin arbitration (same as APB)
                    grant_matrix[s] = '0;
                    for (int i = 0; i < NUM_MASTERS; i++) begin
                        int m;
                        m = (last_grant[s] + 1 + i) % NUM_MASTERS;
                        if (request_matrix[s][m] && grant_matrix[s] == '0) begin
                            grant_matrix[s][m] = 1'b1;
                            last_grant[s] = m[$clog2(NUM_MASTERS)-1:0];
                            packet_active[s] = 1'b1;
                        end
                    end
                end else begin
                    grant_matrix[s] <= '0;
                end
            end
        end
    end
endgenerate

// ==========================================================================
// Crossbar Data Multiplexing
// ==========================================================================
// Same pattern as APB crossbar, just more signals:
// - APB muxes: PRDATA, PSLVERR
// - AXIS muxes: TDATA, TVALID, TLAST, TDEST, TID, TUSER
// ==========================================================================

generate
    for (genvar s = 0; s < NUM_SLAVES; s++) begin : gen_slave_mux
        always_comb begin
            // Default: all zeros
            m_axis_tdata[s]  = '0;
            m_axis_tvalid[s] = 1'b0;
            m_axis_tlast[s]  = 1'b0;
            m_axis_tdest[s]  = '0;
            m_axis_tid[s]    = '0;
            m_axis_tuser[s]  = '0;

            // Multiplex granted master to this slave
            for (int m = 0; m < NUM_MASTERS; m++) begin
                if (grant_matrix[s][m]) begin
                    m_axis_tdata[s]  = s_axis_tdata[m];
                    m_axis_tvalid[s] = s_axis_tvalid[m];
                    m_axis_tlast[s]  = s_axis_tlast[m];
                    m_axis_tdest[s]  = s_axis_tdest[m];
                    m_axis_tid[s]    = s_axis_tid[m];
                    m_axis_tuser[s]  = s_axis_tuser[m];
                end
            end
        end
    end
endgenerate

// ==========================================================================
// Backpressure (TREADY) Logic
// ==========================================================================
// Identical to APB PREADY logic, just renamed signal:
// - APB: pready[m] = pready_slave[granted_slave]
// - AXIS: s_axis_tready[m] = m_axis_tready[granted_slave]
// ==========================================================================

generate
    for (genvar m = 0; m < NUM_MASTERS; m++) begin : gen_master_tready
        always_comb begin
            s_axis_tready[m] = 1'b0;
            for (int s = 0; s < NUM_SLAVES; s++) begin
                if (grant_matrix[s][m]) begin
                    s_axis_tready[m] = m_axis_tready[s];
                end
            end
        end
    end
endgenerate

// ==========================================================================
// Performance Counters (Optional)
// ==========================================================================
// Track packets and transfers per master/slave for performance analysis
// ==========================================================================

// Packet counters per master
logic [31:0] pkt_count_master [NUM_MASTERS];
logic [31:0] pkt_count_slave [NUM_SLAVES];

generate
    // Master packet counters
    for (genvar m = 0; m < NUM_MASTERS; m++) begin : gen_master_counters
        always_ff @(posedge aclk or negedge aresetn) begin
            if (!aresetn)
                pkt_count_master[m] <= '0;
            else if (s_axis_tvalid[m] && s_axis_tready[m] && s_axis_tlast[m])
                pkt_count_master[m] <= pkt_count_master[m] + 1;
        end
    end

    // Slave packet counters
    for (genvar s = 0; s < NUM_SLAVES; s++) begin : gen_slave_counters
        always_ff @(posedge aclk or negedge aresetn) begin
            if (!aresetn)
                pkt_count_slave[s] <= '0;
            else if (m_axis_tvalid[s] && m_axis_tready[s] && m_axis_tlast[s])
                pkt_count_slave[s] <= pkt_count_slave[s] + 1;
        end
    end
endgenerate

// ==========================================================================
// Assertions for Debug and Verification
// ==========================================================================
`ifdef FORMAL
// One-hot grant check
generate
    for (genvar s = 0; s < NUM_SLAVES; s++) begin : gen_onehot_assert
        assert property (@(posedge aclk) disable iff (!aresetn)
            $onehot0(grant_matrix[s])
        ) else $error("Grant matrix not one-hot for slave %0d", s);
    end
endgenerate

// TDEST in range check
generate
    for (genvar m = 0; m < NUM_MASTERS; m++) begin : gen_tdest_assert
        assert property (@(posedge aclk) disable iff (!aresetn)
            s_axis_tvalid[m] |-> s_axis_tdest[m] < NUM_SLAVES
        ) else $error("TDEST out of range for master %0d", m);
    end
endgenerate
`endif

endmodule
