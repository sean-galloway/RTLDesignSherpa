`timescale 1ns / 1ps

// taken from here: https://stackoverflow.com/questions/49527064/sorting-in-verilog-with-one-cycle
// with only minor updates
module sort #(
    parameter NUM_VALS = 5,
    parameter SIZE     = 16
)(  input  logic                     i_clk, i_rst_n,
    input  logic [NUM_VALS*SIZE-1:0] i_data,
    output logic [NUM_VALS*SIZE-1:0] o_data
);
    logic [NUM_VALS*SIZE-1:0] w_sorted_bus;
    always_ff @(posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n)
            o_data <= 'b0;
        else
            o_data <= w_sorted_bus;
    end

    integer i, j;
    logic [SIZE-1:0] w_temp;
    logic [SIZE-1:0] w_array [1:NUM_VALS];
    always_comb begin
        for (i = 0; i < NUM_VALS; i = i + 1) begin
            w_array[i+1] = i_data[i*SIZE +: SIZE];
        end

        for (i = NUM_VALS; i > 0; i = i - 1) begin
            for (j = 1 ; j < i; j = j + 1) begin
                if (w_array[j] < w_array[j + 1]) begin
                    w_temp         = w_array[j];
                    w_array[j]     = w_array[j + 1];
                    w_array[j + 1] = w_temp;
                end 
            end
        end

        for (i = 0; i < NUM_VALS; i = i + 1) begin
            w_sorted_bus[i*SIZE +: SIZE] = w_array[i+1];
        end
    end

    // synopsys translate_off
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, sort);
    end
    // synopsys translate_on
endmodule