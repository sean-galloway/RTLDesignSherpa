`timescale 1ns / 1ps

module math_adder_brent_kung_grouppg_008 #(parameter   N = 8)(
    input  logic [N:0] i_p,
    input  logic [N:0] i_g,
    output logic [N:0] ow_gg,
    output logic [N:0] ow_pp
);

logic  G_3_2;
logic  P_3_2;
logic  G_5_4;
logic  P_5_4;
logic  G_7_6;
logic  P_7_6;
logic  G_7_4;
logic  P_7_4;
math_adder_brent_kung_gray gray_block_1_0(.i_g(i_g[1]),.i_p(i_p[1]),.i_g_km1(i_g[0]),.ow_g(ow_gg[1]));
math_adder_brent_kung_black black_block_3_2(.i_g(i_g[3]),.i_p(i_p[3]),.i_g_km1(i_g[2]),.i_p_km1(i_p[2]),.ow_g(G_3_2),.ow_p(P_3_2));
math_adder_brent_kung_black black_block_5_4(.i_g(i_g[5]),.i_p(i_p[5]),.i_g_km1(i_g[4]),.i_p_km1(i_p[4]),.ow_g(G_5_4),.ow_p(P_5_4));
math_adder_brent_kung_black black_block_7_6(.i_g(i_g[7]),.i_p(i_p[7]),.i_g_km1(i_g[6]),.i_p_km1(i_p[6]),.ow_g(G_7_6),.ow_p(P_7_6));
math_adder_brent_kung_gray gray_block_3_0(.i_g(G_3_2),.i_p(P_3_2),.i_g_km1(ow_gg[1]),.ow_g(ow_gg[3]));
math_adder_brent_kung_black black_block_7_4(.i_g(G_7_6),.i_p(P_7_6),.i_g_km1(G_5_4),.i_p_km1(P_5_4),.ow_g(G_7_4),.ow_p(P_7_4));
math_adder_brent_kung_gray gray_block_7_0(.i_g(G_7_4),.i_p(P_7_4),.i_g_km1(ow_gg[3]),.ow_g(ow_gg[7]));
math_adder_brent_kung_gray gray_block_5_3(.i_g(G_5_4),.i_p(P_5_4),.i_g_km1(ow_gg[3]),.ow_g(ow_gg[5]));
math_adder_brent_kung_gray gray_block_2_1(.i_g(i_g[2]),.i_p(i_p[2]),.i_g_km1(ow_gg[1]),.ow_g(ow_gg[2]));
math_adder_brent_kung_gray gray_block_4_3(.i_g(i_g[4]),.i_p(i_p[4]),.i_g_km1(ow_gg[3]),.ow_g(ow_gg[4]));
math_adder_brent_kung_gray gray_block_6_5(.i_g(i_g[6]),.i_p(i_p[6]),.i_g_km1(ow_gg[5]),.ow_g(ow_gg[6]));
math_adder_brent_kung_gray gray_block_8_7(.i_g(i_g[8]),.i_p(i_p[8]),.i_g_km1(ow_gg[7]),.ow_g(ow_gg[8]));
assign ow_gg[0] = i_g[0];
assign ow_pp[0] = i_p[0];
endmodule
