../amba/includes/monitor_pkg.sv