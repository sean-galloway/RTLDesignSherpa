`timescale 1ns / 1ps

module math_multiplier_wallace_tree_032 (
    input  [31:0] i_multiplier,
    input  [31:0] i_multiplicand,
    output [63:0] ow_product
);

// Partial products generation
wire w_pp_00_00 = i_multiplier[ 0] & i_multiplicand[ 0];
wire w_pp_00_01 = i_multiplier[ 0] & i_multiplicand[ 1];
wire w_pp_00_02 = i_multiplier[ 0] & i_multiplicand[ 2];
wire w_pp_00_03 = i_multiplier[ 0] & i_multiplicand[ 3];
wire w_pp_00_04 = i_multiplier[ 0] & i_multiplicand[ 4];
wire w_pp_00_05 = i_multiplier[ 0] & i_multiplicand[ 5];
wire w_pp_00_06 = i_multiplier[ 0] & i_multiplicand[ 6];
wire w_pp_00_07 = i_multiplier[ 0] & i_multiplicand[ 7];
wire w_pp_00_08 = i_multiplier[ 0] & i_multiplicand[ 8];
wire w_pp_00_09 = i_multiplier[ 0] & i_multiplicand[ 9];
wire w_pp_00_10 = i_multiplier[ 0] & i_multiplicand[10];
wire w_pp_00_11 = i_multiplier[ 0] & i_multiplicand[11];
wire w_pp_00_12 = i_multiplier[ 0] & i_multiplicand[12];
wire w_pp_00_13 = i_multiplier[ 0] & i_multiplicand[13];
wire w_pp_00_14 = i_multiplier[ 0] & i_multiplicand[14];
wire w_pp_00_15 = i_multiplier[ 0] & i_multiplicand[15];
wire w_pp_00_16 = i_multiplier[ 0] & i_multiplicand[16];
wire w_pp_00_17 = i_multiplier[ 0] & i_multiplicand[17];
wire w_pp_00_18 = i_multiplier[ 0] & i_multiplicand[18];
wire w_pp_00_19 = i_multiplier[ 0] & i_multiplicand[19];
wire w_pp_00_20 = i_multiplier[ 0] & i_multiplicand[20];
wire w_pp_00_21 = i_multiplier[ 0] & i_multiplicand[21];
wire w_pp_00_22 = i_multiplier[ 0] & i_multiplicand[22];
wire w_pp_00_23 = i_multiplier[ 0] & i_multiplicand[23];
wire w_pp_00_24 = i_multiplier[ 0] & i_multiplicand[24];
wire w_pp_00_25 = i_multiplier[ 0] & i_multiplicand[25];
wire w_pp_00_26 = i_multiplier[ 0] & i_multiplicand[26];
wire w_pp_00_27 = i_multiplier[ 0] & i_multiplicand[27];
wire w_pp_00_28 = i_multiplier[ 0] & i_multiplicand[28];
wire w_pp_00_29 = i_multiplier[ 0] & i_multiplicand[29];
wire w_pp_00_30 = i_multiplier[ 0] & i_multiplicand[30];
wire w_pp_00_31 = i_multiplier[ 0] & i_multiplicand[31];
wire w_pp_01_00 = i_multiplier[ 1] & i_multiplicand[ 0];
wire w_pp_01_01 = i_multiplier[ 1] & i_multiplicand[ 1];
wire w_pp_01_02 = i_multiplier[ 1] & i_multiplicand[ 2];
wire w_pp_01_03 = i_multiplier[ 1] & i_multiplicand[ 3];
wire w_pp_01_04 = i_multiplier[ 1] & i_multiplicand[ 4];
wire w_pp_01_05 = i_multiplier[ 1] & i_multiplicand[ 5];
wire w_pp_01_06 = i_multiplier[ 1] & i_multiplicand[ 6];
wire w_pp_01_07 = i_multiplier[ 1] & i_multiplicand[ 7];
wire w_pp_01_08 = i_multiplier[ 1] & i_multiplicand[ 8];
wire w_pp_01_09 = i_multiplier[ 1] & i_multiplicand[ 9];
wire w_pp_01_10 = i_multiplier[ 1] & i_multiplicand[10];
wire w_pp_01_11 = i_multiplier[ 1] & i_multiplicand[11];
wire w_pp_01_12 = i_multiplier[ 1] & i_multiplicand[12];
wire w_pp_01_13 = i_multiplier[ 1] & i_multiplicand[13];
wire w_pp_01_14 = i_multiplier[ 1] & i_multiplicand[14];
wire w_pp_01_15 = i_multiplier[ 1] & i_multiplicand[15];
wire w_pp_01_16 = i_multiplier[ 1] & i_multiplicand[16];
wire w_pp_01_17 = i_multiplier[ 1] & i_multiplicand[17];
wire w_pp_01_18 = i_multiplier[ 1] & i_multiplicand[18];
wire w_pp_01_19 = i_multiplier[ 1] & i_multiplicand[19];
wire w_pp_01_20 = i_multiplier[ 1] & i_multiplicand[20];
wire w_pp_01_21 = i_multiplier[ 1] & i_multiplicand[21];
wire w_pp_01_22 = i_multiplier[ 1] & i_multiplicand[22];
wire w_pp_01_23 = i_multiplier[ 1] & i_multiplicand[23];
wire w_pp_01_24 = i_multiplier[ 1] & i_multiplicand[24];
wire w_pp_01_25 = i_multiplier[ 1] & i_multiplicand[25];
wire w_pp_01_26 = i_multiplier[ 1] & i_multiplicand[26];
wire w_pp_01_27 = i_multiplier[ 1] & i_multiplicand[27];
wire w_pp_01_28 = i_multiplier[ 1] & i_multiplicand[28];
wire w_pp_01_29 = i_multiplier[ 1] & i_multiplicand[29];
wire w_pp_01_30 = i_multiplier[ 1] & i_multiplicand[30];
wire w_pp_01_31 = i_multiplier[ 1] & i_multiplicand[31];
wire w_pp_02_00 = i_multiplier[ 2] & i_multiplicand[ 0];
wire w_pp_02_01 = i_multiplier[ 2] & i_multiplicand[ 1];
wire w_pp_02_02 = i_multiplier[ 2] & i_multiplicand[ 2];
wire w_pp_02_03 = i_multiplier[ 2] & i_multiplicand[ 3];
wire w_pp_02_04 = i_multiplier[ 2] & i_multiplicand[ 4];
wire w_pp_02_05 = i_multiplier[ 2] & i_multiplicand[ 5];
wire w_pp_02_06 = i_multiplier[ 2] & i_multiplicand[ 6];
wire w_pp_02_07 = i_multiplier[ 2] & i_multiplicand[ 7];
wire w_pp_02_08 = i_multiplier[ 2] & i_multiplicand[ 8];
wire w_pp_02_09 = i_multiplier[ 2] & i_multiplicand[ 9];
wire w_pp_02_10 = i_multiplier[ 2] & i_multiplicand[10];
wire w_pp_02_11 = i_multiplier[ 2] & i_multiplicand[11];
wire w_pp_02_12 = i_multiplier[ 2] & i_multiplicand[12];
wire w_pp_02_13 = i_multiplier[ 2] & i_multiplicand[13];
wire w_pp_02_14 = i_multiplier[ 2] & i_multiplicand[14];
wire w_pp_02_15 = i_multiplier[ 2] & i_multiplicand[15];
wire w_pp_02_16 = i_multiplier[ 2] & i_multiplicand[16];
wire w_pp_02_17 = i_multiplier[ 2] & i_multiplicand[17];
wire w_pp_02_18 = i_multiplier[ 2] & i_multiplicand[18];
wire w_pp_02_19 = i_multiplier[ 2] & i_multiplicand[19];
wire w_pp_02_20 = i_multiplier[ 2] & i_multiplicand[20];
wire w_pp_02_21 = i_multiplier[ 2] & i_multiplicand[21];
wire w_pp_02_22 = i_multiplier[ 2] & i_multiplicand[22];
wire w_pp_02_23 = i_multiplier[ 2] & i_multiplicand[23];
wire w_pp_02_24 = i_multiplier[ 2] & i_multiplicand[24];
wire w_pp_02_25 = i_multiplier[ 2] & i_multiplicand[25];
wire w_pp_02_26 = i_multiplier[ 2] & i_multiplicand[26];
wire w_pp_02_27 = i_multiplier[ 2] & i_multiplicand[27];
wire w_pp_02_28 = i_multiplier[ 2] & i_multiplicand[28];
wire w_pp_02_29 = i_multiplier[ 2] & i_multiplicand[29];
wire w_pp_02_30 = i_multiplier[ 2] & i_multiplicand[30];
wire w_pp_02_31 = i_multiplier[ 2] & i_multiplicand[31];
wire w_pp_03_00 = i_multiplier[ 3] & i_multiplicand[ 0];
wire w_pp_03_01 = i_multiplier[ 3] & i_multiplicand[ 1];
wire w_pp_03_02 = i_multiplier[ 3] & i_multiplicand[ 2];
wire w_pp_03_03 = i_multiplier[ 3] & i_multiplicand[ 3];
wire w_pp_03_04 = i_multiplier[ 3] & i_multiplicand[ 4];
wire w_pp_03_05 = i_multiplier[ 3] & i_multiplicand[ 5];
wire w_pp_03_06 = i_multiplier[ 3] & i_multiplicand[ 6];
wire w_pp_03_07 = i_multiplier[ 3] & i_multiplicand[ 7];
wire w_pp_03_08 = i_multiplier[ 3] & i_multiplicand[ 8];
wire w_pp_03_09 = i_multiplier[ 3] & i_multiplicand[ 9];
wire w_pp_03_10 = i_multiplier[ 3] & i_multiplicand[10];
wire w_pp_03_11 = i_multiplier[ 3] & i_multiplicand[11];
wire w_pp_03_12 = i_multiplier[ 3] & i_multiplicand[12];
wire w_pp_03_13 = i_multiplier[ 3] & i_multiplicand[13];
wire w_pp_03_14 = i_multiplier[ 3] & i_multiplicand[14];
wire w_pp_03_15 = i_multiplier[ 3] & i_multiplicand[15];
wire w_pp_03_16 = i_multiplier[ 3] & i_multiplicand[16];
wire w_pp_03_17 = i_multiplier[ 3] & i_multiplicand[17];
wire w_pp_03_18 = i_multiplier[ 3] & i_multiplicand[18];
wire w_pp_03_19 = i_multiplier[ 3] & i_multiplicand[19];
wire w_pp_03_20 = i_multiplier[ 3] & i_multiplicand[20];
wire w_pp_03_21 = i_multiplier[ 3] & i_multiplicand[21];
wire w_pp_03_22 = i_multiplier[ 3] & i_multiplicand[22];
wire w_pp_03_23 = i_multiplier[ 3] & i_multiplicand[23];
wire w_pp_03_24 = i_multiplier[ 3] & i_multiplicand[24];
wire w_pp_03_25 = i_multiplier[ 3] & i_multiplicand[25];
wire w_pp_03_26 = i_multiplier[ 3] & i_multiplicand[26];
wire w_pp_03_27 = i_multiplier[ 3] & i_multiplicand[27];
wire w_pp_03_28 = i_multiplier[ 3] & i_multiplicand[28];
wire w_pp_03_29 = i_multiplier[ 3] & i_multiplicand[29];
wire w_pp_03_30 = i_multiplier[ 3] & i_multiplicand[30];
wire w_pp_03_31 = i_multiplier[ 3] & i_multiplicand[31];
wire w_pp_04_00 = i_multiplier[ 4] & i_multiplicand[ 0];
wire w_pp_04_01 = i_multiplier[ 4] & i_multiplicand[ 1];
wire w_pp_04_02 = i_multiplier[ 4] & i_multiplicand[ 2];
wire w_pp_04_03 = i_multiplier[ 4] & i_multiplicand[ 3];
wire w_pp_04_04 = i_multiplier[ 4] & i_multiplicand[ 4];
wire w_pp_04_05 = i_multiplier[ 4] & i_multiplicand[ 5];
wire w_pp_04_06 = i_multiplier[ 4] & i_multiplicand[ 6];
wire w_pp_04_07 = i_multiplier[ 4] & i_multiplicand[ 7];
wire w_pp_04_08 = i_multiplier[ 4] & i_multiplicand[ 8];
wire w_pp_04_09 = i_multiplier[ 4] & i_multiplicand[ 9];
wire w_pp_04_10 = i_multiplier[ 4] & i_multiplicand[10];
wire w_pp_04_11 = i_multiplier[ 4] & i_multiplicand[11];
wire w_pp_04_12 = i_multiplier[ 4] & i_multiplicand[12];
wire w_pp_04_13 = i_multiplier[ 4] & i_multiplicand[13];
wire w_pp_04_14 = i_multiplier[ 4] & i_multiplicand[14];
wire w_pp_04_15 = i_multiplier[ 4] & i_multiplicand[15];
wire w_pp_04_16 = i_multiplier[ 4] & i_multiplicand[16];
wire w_pp_04_17 = i_multiplier[ 4] & i_multiplicand[17];
wire w_pp_04_18 = i_multiplier[ 4] & i_multiplicand[18];
wire w_pp_04_19 = i_multiplier[ 4] & i_multiplicand[19];
wire w_pp_04_20 = i_multiplier[ 4] & i_multiplicand[20];
wire w_pp_04_21 = i_multiplier[ 4] & i_multiplicand[21];
wire w_pp_04_22 = i_multiplier[ 4] & i_multiplicand[22];
wire w_pp_04_23 = i_multiplier[ 4] & i_multiplicand[23];
wire w_pp_04_24 = i_multiplier[ 4] & i_multiplicand[24];
wire w_pp_04_25 = i_multiplier[ 4] & i_multiplicand[25];
wire w_pp_04_26 = i_multiplier[ 4] & i_multiplicand[26];
wire w_pp_04_27 = i_multiplier[ 4] & i_multiplicand[27];
wire w_pp_04_28 = i_multiplier[ 4] & i_multiplicand[28];
wire w_pp_04_29 = i_multiplier[ 4] & i_multiplicand[29];
wire w_pp_04_30 = i_multiplier[ 4] & i_multiplicand[30];
wire w_pp_04_31 = i_multiplier[ 4] & i_multiplicand[31];
wire w_pp_05_00 = i_multiplier[ 5] & i_multiplicand[ 0];
wire w_pp_05_01 = i_multiplier[ 5] & i_multiplicand[ 1];
wire w_pp_05_02 = i_multiplier[ 5] & i_multiplicand[ 2];
wire w_pp_05_03 = i_multiplier[ 5] & i_multiplicand[ 3];
wire w_pp_05_04 = i_multiplier[ 5] & i_multiplicand[ 4];
wire w_pp_05_05 = i_multiplier[ 5] & i_multiplicand[ 5];
wire w_pp_05_06 = i_multiplier[ 5] & i_multiplicand[ 6];
wire w_pp_05_07 = i_multiplier[ 5] & i_multiplicand[ 7];
wire w_pp_05_08 = i_multiplier[ 5] & i_multiplicand[ 8];
wire w_pp_05_09 = i_multiplier[ 5] & i_multiplicand[ 9];
wire w_pp_05_10 = i_multiplier[ 5] & i_multiplicand[10];
wire w_pp_05_11 = i_multiplier[ 5] & i_multiplicand[11];
wire w_pp_05_12 = i_multiplier[ 5] & i_multiplicand[12];
wire w_pp_05_13 = i_multiplier[ 5] & i_multiplicand[13];
wire w_pp_05_14 = i_multiplier[ 5] & i_multiplicand[14];
wire w_pp_05_15 = i_multiplier[ 5] & i_multiplicand[15];
wire w_pp_05_16 = i_multiplier[ 5] & i_multiplicand[16];
wire w_pp_05_17 = i_multiplier[ 5] & i_multiplicand[17];
wire w_pp_05_18 = i_multiplier[ 5] & i_multiplicand[18];
wire w_pp_05_19 = i_multiplier[ 5] & i_multiplicand[19];
wire w_pp_05_20 = i_multiplier[ 5] & i_multiplicand[20];
wire w_pp_05_21 = i_multiplier[ 5] & i_multiplicand[21];
wire w_pp_05_22 = i_multiplier[ 5] & i_multiplicand[22];
wire w_pp_05_23 = i_multiplier[ 5] & i_multiplicand[23];
wire w_pp_05_24 = i_multiplier[ 5] & i_multiplicand[24];
wire w_pp_05_25 = i_multiplier[ 5] & i_multiplicand[25];
wire w_pp_05_26 = i_multiplier[ 5] & i_multiplicand[26];
wire w_pp_05_27 = i_multiplier[ 5] & i_multiplicand[27];
wire w_pp_05_28 = i_multiplier[ 5] & i_multiplicand[28];
wire w_pp_05_29 = i_multiplier[ 5] & i_multiplicand[29];
wire w_pp_05_30 = i_multiplier[ 5] & i_multiplicand[30];
wire w_pp_05_31 = i_multiplier[ 5] & i_multiplicand[31];
wire w_pp_06_00 = i_multiplier[ 6] & i_multiplicand[ 0];
wire w_pp_06_01 = i_multiplier[ 6] & i_multiplicand[ 1];
wire w_pp_06_02 = i_multiplier[ 6] & i_multiplicand[ 2];
wire w_pp_06_03 = i_multiplier[ 6] & i_multiplicand[ 3];
wire w_pp_06_04 = i_multiplier[ 6] & i_multiplicand[ 4];
wire w_pp_06_05 = i_multiplier[ 6] & i_multiplicand[ 5];
wire w_pp_06_06 = i_multiplier[ 6] & i_multiplicand[ 6];
wire w_pp_06_07 = i_multiplier[ 6] & i_multiplicand[ 7];
wire w_pp_06_08 = i_multiplier[ 6] & i_multiplicand[ 8];
wire w_pp_06_09 = i_multiplier[ 6] & i_multiplicand[ 9];
wire w_pp_06_10 = i_multiplier[ 6] & i_multiplicand[10];
wire w_pp_06_11 = i_multiplier[ 6] & i_multiplicand[11];
wire w_pp_06_12 = i_multiplier[ 6] & i_multiplicand[12];
wire w_pp_06_13 = i_multiplier[ 6] & i_multiplicand[13];
wire w_pp_06_14 = i_multiplier[ 6] & i_multiplicand[14];
wire w_pp_06_15 = i_multiplier[ 6] & i_multiplicand[15];
wire w_pp_06_16 = i_multiplier[ 6] & i_multiplicand[16];
wire w_pp_06_17 = i_multiplier[ 6] & i_multiplicand[17];
wire w_pp_06_18 = i_multiplier[ 6] & i_multiplicand[18];
wire w_pp_06_19 = i_multiplier[ 6] & i_multiplicand[19];
wire w_pp_06_20 = i_multiplier[ 6] & i_multiplicand[20];
wire w_pp_06_21 = i_multiplier[ 6] & i_multiplicand[21];
wire w_pp_06_22 = i_multiplier[ 6] & i_multiplicand[22];
wire w_pp_06_23 = i_multiplier[ 6] & i_multiplicand[23];
wire w_pp_06_24 = i_multiplier[ 6] & i_multiplicand[24];
wire w_pp_06_25 = i_multiplier[ 6] & i_multiplicand[25];
wire w_pp_06_26 = i_multiplier[ 6] & i_multiplicand[26];
wire w_pp_06_27 = i_multiplier[ 6] & i_multiplicand[27];
wire w_pp_06_28 = i_multiplier[ 6] & i_multiplicand[28];
wire w_pp_06_29 = i_multiplier[ 6] & i_multiplicand[29];
wire w_pp_06_30 = i_multiplier[ 6] & i_multiplicand[30];
wire w_pp_06_31 = i_multiplier[ 6] & i_multiplicand[31];
wire w_pp_07_00 = i_multiplier[ 7] & i_multiplicand[ 0];
wire w_pp_07_01 = i_multiplier[ 7] & i_multiplicand[ 1];
wire w_pp_07_02 = i_multiplier[ 7] & i_multiplicand[ 2];
wire w_pp_07_03 = i_multiplier[ 7] & i_multiplicand[ 3];
wire w_pp_07_04 = i_multiplier[ 7] & i_multiplicand[ 4];
wire w_pp_07_05 = i_multiplier[ 7] & i_multiplicand[ 5];
wire w_pp_07_06 = i_multiplier[ 7] & i_multiplicand[ 6];
wire w_pp_07_07 = i_multiplier[ 7] & i_multiplicand[ 7];
wire w_pp_07_08 = i_multiplier[ 7] & i_multiplicand[ 8];
wire w_pp_07_09 = i_multiplier[ 7] & i_multiplicand[ 9];
wire w_pp_07_10 = i_multiplier[ 7] & i_multiplicand[10];
wire w_pp_07_11 = i_multiplier[ 7] & i_multiplicand[11];
wire w_pp_07_12 = i_multiplier[ 7] & i_multiplicand[12];
wire w_pp_07_13 = i_multiplier[ 7] & i_multiplicand[13];
wire w_pp_07_14 = i_multiplier[ 7] & i_multiplicand[14];
wire w_pp_07_15 = i_multiplier[ 7] & i_multiplicand[15];
wire w_pp_07_16 = i_multiplier[ 7] & i_multiplicand[16];
wire w_pp_07_17 = i_multiplier[ 7] & i_multiplicand[17];
wire w_pp_07_18 = i_multiplier[ 7] & i_multiplicand[18];
wire w_pp_07_19 = i_multiplier[ 7] & i_multiplicand[19];
wire w_pp_07_20 = i_multiplier[ 7] & i_multiplicand[20];
wire w_pp_07_21 = i_multiplier[ 7] & i_multiplicand[21];
wire w_pp_07_22 = i_multiplier[ 7] & i_multiplicand[22];
wire w_pp_07_23 = i_multiplier[ 7] & i_multiplicand[23];
wire w_pp_07_24 = i_multiplier[ 7] & i_multiplicand[24];
wire w_pp_07_25 = i_multiplier[ 7] & i_multiplicand[25];
wire w_pp_07_26 = i_multiplier[ 7] & i_multiplicand[26];
wire w_pp_07_27 = i_multiplier[ 7] & i_multiplicand[27];
wire w_pp_07_28 = i_multiplier[ 7] & i_multiplicand[28];
wire w_pp_07_29 = i_multiplier[ 7] & i_multiplicand[29];
wire w_pp_07_30 = i_multiplier[ 7] & i_multiplicand[30];
wire w_pp_07_31 = i_multiplier[ 7] & i_multiplicand[31];
wire w_pp_08_00 = i_multiplier[ 8] & i_multiplicand[ 0];
wire w_pp_08_01 = i_multiplier[ 8] & i_multiplicand[ 1];
wire w_pp_08_02 = i_multiplier[ 8] & i_multiplicand[ 2];
wire w_pp_08_03 = i_multiplier[ 8] & i_multiplicand[ 3];
wire w_pp_08_04 = i_multiplier[ 8] & i_multiplicand[ 4];
wire w_pp_08_05 = i_multiplier[ 8] & i_multiplicand[ 5];
wire w_pp_08_06 = i_multiplier[ 8] & i_multiplicand[ 6];
wire w_pp_08_07 = i_multiplier[ 8] & i_multiplicand[ 7];
wire w_pp_08_08 = i_multiplier[ 8] & i_multiplicand[ 8];
wire w_pp_08_09 = i_multiplier[ 8] & i_multiplicand[ 9];
wire w_pp_08_10 = i_multiplier[ 8] & i_multiplicand[10];
wire w_pp_08_11 = i_multiplier[ 8] & i_multiplicand[11];
wire w_pp_08_12 = i_multiplier[ 8] & i_multiplicand[12];
wire w_pp_08_13 = i_multiplier[ 8] & i_multiplicand[13];
wire w_pp_08_14 = i_multiplier[ 8] & i_multiplicand[14];
wire w_pp_08_15 = i_multiplier[ 8] & i_multiplicand[15];
wire w_pp_08_16 = i_multiplier[ 8] & i_multiplicand[16];
wire w_pp_08_17 = i_multiplier[ 8] & i_multiplicand[17];
wire w_pp_08_18 = i_multiplier[ 8] & i_multiplicand[18];
wire w_pp_08_19 = i_multiplier[ 8] & i_multiplicand[19];
wire w_pp_08_20 = i_multiplier[ 8] & i_multiplicand[20];
wire w_pp_08_21 = i_multiplier[ 8] & i_multiplicand[21];
wire w_pp_08_22 = i_multiplier[ 8] & i_multiplicand[22];
wire w_pp_08_23 = i_multiplier[ 8] & i_multiplicand[23];
wire w_pp_08_24 = i_multiplier[ 8] & i_multiplicand[24];
wire w_pp_08_25 = i_multiplier[ 8] & i_multiplicand[25];
wire w_pp_08_26 = i_multiplier[ 8] & i_multiplicand[26];
wire w_pp_08_27 = i_multiplier[ 8] & i_multiplicand[27];
wire w_pp_08_28 = i_multiplier[ 8] & i_multiplicand[28];
wire w_pp_08_29 = i_multiplier[ 8] & i_multiplicand[29];
wire w_pp_08_30 = i_multiplier[ 8] & i_multiplicand[30];
wire w_pp_08_31 = i_multiplier[ 8] & i_multiplicand[31];
wire w_pp_09_00 = i_multiplier[ 9] & i_multiplicand[ 0];
wire w_pp_09_01 = i_multiplier[ 9] & i_multiplicand[ 1];
wire w_pp_09_02 = i_multiplier[ 9] & i_multiplicand[ 2];
wire w_pp_09_03 = i_multiplier[ 9] & i_multiplicand[ 3];
wire w_pp_09_04 = i_multiplier[ 9] & i_multiplicand[ 4];
wire w_pp_09_05 = i_multiplier[ 9] & i_multiplicand[ 5];
wire w_pp_09_06 = i_multiplier[ 9] & i_multiplicand[ 6];
wire w_pp_09_07 = i_multiplier[ 9] & i_multiplicand[ 7];
wire w_pp_09_08 = i_multiplier[ 9] & i_multiplicand[ 8];
wire w_pp_09_09 = i_multiplier[ 9] & i_multiplicand[ 9];
wire w_pp_09_10 = i_multiplier[ 9] & i_multiplicand[10];
wire w_pp_09_11 = i_multiplier[ 9] & i_multiplicand[11];
wire w_pp_09_12 = i_multiplier[ 9] & i_multiplicand[12];
wire w_pp_09_13 = i_multiplier[ 9] & i_multiplicand[13];
wire w_pp_09_14 = i_multiplier[ 9] & i_multiplicand[14];
wire w_pp_09_15 = i_multiplier[ 9] & i_multiplicand[15];
wire w_pp_09_16 = i_multiplier[ 9] & i_multiplicand[16];
wire w_pp_09_17 = i_multiplier[ 9] & i_multiplicand[17];
wire w_pp_09_18 = i_multiplier[ 9] & i_multiplicand[18];
wire w_pp_09_19 = i_multiplier[ 9] & i_multiplicand[19];
wire w_pp_09_20 = i_multiplier[ 9] & i_multiplicand[20];
wire w_pp_09_21 = i_multiplier[ 9] & i_multiplicand[21];
wire w_pp_09_22 = i_multiplier[ 9] & i_multiplicand[22];
wire w_pp_09_23 = i_multiplier[ 9] & i_multiplicand[23];
wire w_pp_09_24 = i_multiplier[ 9] & i_multiplicand[24];
wire w_pp_09_25 = i_multiplier[ 9] & i_multiplicand[25];
wire w_pp_09_26 = i_multiplier[ 9] & i_multiplicand[26];
wire w_pp_09_27 = i_multiplier[ 9] & i_multiplicand[27];
wire w_pp_09_28 = i_multiplier[ 9] & i_multiplicand[28];
wire w_pp_09_29 = i_multiplier[ 9] & i_multiplicand[29];
wire w_pp_09_30 = i_multiplier[ 9] & i_multiplicand[30];
wire w_pp_09_31 = i_multiplier[ 9] & i_multiplicand[31];
wire w_pp_10_00 = i_multiplier[10] & i_multiplicand[ 0];
wire w_pp_10_01 = i_multiplier[10] & i_multiplicand[ 1];
wire w_pp_10_02 = i_multiplier[10] & i_multiplicand[ 2];
wire w_pp_10_03 = i_multiplier[10] & i_multiplicand[ 3];
wire w_pp_10_04 = i_multiplier[10] & i_multiplicand[ 4];
wire w_pp_10_05 = i_multiplier[10] & i_multiplicand[ 5];
wire w_pp_10_06 = i_multiplier[10] & i_multiplicand[ 6];
wire w_pp_10_07 = i_multiplier[10] & i_multiplicand[ 7];
wire w_pp_10_08 = i_multiplier[10] & i_multiplicand[ 8];
wire w_pp_10_09 = i_multiplier[10] & i_multiplicand[ 9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_10_16 = i_multiplier[10] & i_multiplicand[16];
wire w_pp_10_17 = i_multiplier[10] & i_multiplicand[17];
wire w_pp_10_18 = i_multiplier[10] & i_multiplicand[18];
wire w_pp_10_19 = i_multiplier[10] & i_multiplicand[19];
wire w_pp_10_20 = i_multiplier[10] & i_multiplicand[20];
wire w_pp_10_21 = i_multiplier[10] & i_multiplicand[21];
wire w_pp_10_22 = i_multiplier[10] & i_multiplicand[22];
wire w_pp_10_23 = i_multiplier[10] & i_multiplicand[23];
wire w_pp_10_24 = i_multiplier[10] & i_multiplicand[24];
wire w_pp_10_25 = i_multiplier[10] & i_multiplicand[25];
wire w_pp_10_26 = i_multiplier[10] & i_multiplicand[26];
wire w_pp_10_27 = i_multiplier[10] & i_multiplicand[27];
wire w_pp_10_28 = i_multiplier[10] & i_multiplicand[28];
wire w_pp_10_29 = i_multiplier[10] & i_multiplicand[29];
wire w_pp_10_30 = i_multiplier[10] & i_multiplicand[30];
wire w_pp_10_31 = i_multiplier[10] & i_multiplicand[31];
wire w_pp_11_00 = i_multiplier[11] & i_multiplicand[ 0];
wire w_pp_11_01 = i_multiplier[11] & i_multiplicand[ 1];
wire w_pp_11_02 = i_multiplier[11] & i_multiplicand[ 2];
wire w_pp_11_03 = i_multiplier[11] & i_multiplicand[ 3];
wire w_pp_11_04 = i_multiplier[11] & i_multiplicand[ 4];
wire w_pp_11_05 = i_multiplier[11] & i_multiplicand[ 5];
wire w_pp_11_06 = i_multiplier[11] & i_multiplicand[ 6];
wire w_pp_11_07 = i_multiplier[11] & i_multiplicand[ 7];
wire w_pp_11_08 = i_multiplier[11] & i_multiplicand[ 8];
wire w_pp_11_09 = i_multiplier[11] & i_multiplicand[ 9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_11_16 = i_multiplier[11] & i_multiplicand[16];
wire w_pp_11_17 = i_multiplier[11] & i_multiplicand[17];
wire w_pp_11_18 = i_multiplier[11] & i_multiplicand[18];
wire w_pp_11_19 = i_multiplier[11] & i_multiplicand[19];
wire w_pp_11_20 = i_multiplier[11] & i_multiplicand[20];
wire w_pp_11_21 = i_multiplier[11] & i_multiplicand[21];
wire w_pp_11_22 = i_multiplier[11] & i_multiplicand[22];
wire w_pp_11_23 = i_multiplier[11] & i_multiplicand[23];
wire w_pp_11_24 = i_multiplier[11] & i_multiplicand[24];
wire w_pp_11_25 = i_multiplier[11] & i_multiplicand[25];
wire w_pp_11_26 = i_multiplier[11] & i_multiplicand[26];
wire w_pp_11_27 = i_multiplier[11] & i_multiplicand[27];
wire w_pp_11_28 = i_multiplier[11] & i_multiplicand[28];
wire w_pp_11_29 = i_multiplier[11] & i_multiplicand[29];
wire w_pp_11_30 = i_multiplier[11] & i_multiplicand[30];
wire w_pp_11_31 = i_multiplier[11] & i_multiplicand[31];
wire w_pp_12_00 = i_multiplier[12] & i_multiplicand[ 0];
wire w_pp_12_01 = i_multiplier[12] & i_multiplicand[ 1];
wire w_pp_12_02 = i_multiplier[12] & i_multiplicand[ 2];
wire w_pp_12_03 = i_multiplier[12] & i_multiplicand[ 3];
wire w_pp_12_04 = i_multiplier[12] & i_multiplicand[ 4];
wire w_pp_12_05 = i_multiplier[12] & i_multiplicand[ 5];
wire w_pp_12_06 = i_multiplier[12] & i_multiplicand[ 6];
wire w_pp_12_07 = i_multiplier[12] & i_multiplicand[ 7];
wire w_pp_12_08 = i_multiplier[12] & i_multiplicand[ 8];
wire w_pp_12_09 = i_multiplier[12] & i_multiplicand[ 9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_12_16 = i_multiplier[12] & i_multiplicand[16];
wire w_pp_12_17 = i_multiplier[12] & i_multiplicand[17];
wire w_pp_12_18 = i_multiplier[12] & i_multiplicand[18];
wire w_pp_12_19 = i_multiplier[12] & i_multiplicand[19];
wire w_pp_12_20 = i_multiplier[12] & i_multiplicand[20];
wire w_pp_12_21 = i_multiplier[12] & i_multiplicand[21];
wire w_pp_12_22 = i_multiplier[12] & i_multiplicand[22];
wire w_pp_12_23 = i_multiplier[12] & i_multiplicand[23];
wire w_pp_12_24 = i_multiplier[12] & i_multiplicand[24];
wire w_pp_12_25 = i_multiplier[12] & i_multiplicand[25];
wire w_pp_12_26 = i_multiplier[12] & i_multiplicand[26];
wire w_pp_12_27 = i_multiplier[12] & i_multiplicand[27];
wire w_pp_12_28 = i_multiplier[12] & i_multiplicand[28];
wire w_pp_12_29 = i_multiplier[12] & i_multiplicand[29];
wire w_pp_12_30 = i_multiplier[12] & i_multiplicand[30];
wire w_pp_12_31 = i_multiplier[12] & i_multiplicand[31];
wire w_pp_13_00 = i_multiplier[13] & i_multiplicand[ 0];
wire w_pp_13_01 = i_multiplier[13] & i_multiplicand[ 1];
wire w_pp_13_02 = i_multiplier[13] & i_multiplicand[ 2];
wire w_pp_13_03 = i_multiplier[13] & i_multiplicand[ 3];
wire w_pp_13_04 = i_multiplier[13] & i_multiplicand[ 4];
wire w_pp_13_05 = i_multiplier[13] & i_multiplicand[ 5];
wire w_pp_13_06 = i_multiplier[13] & i_multiplicand[ 6];
wire w_pp_13_07 = i_multiplier[13] & i_multiplicand[ 7];
wire w_pp_13_08 = i_multiplier[13] & i_multiplicand[ 8];
wire w_pp_13_09 = i_multiplier[13] & i_multiplicand[ 9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_13_16 = i_multiplier[13] & i_multiplicand[16];
wire w_pp_13_17 = i_multiplier[13] & i_multiplicand[17];
wire w_pp_13_18 = i_multiplier[13] & i_multiplicand[18];
wire w_pp_13_19 = i_multiplier[13] & i_multiplicand[19];
wire w_pp_13_20 = i_multiplier[13] & i_multiplicand[20];
wire w_pp_13_21 = i_multiplier[13] & i_multiplicand[21];
wire w_pp_13_22 = i_multiplier[13] & i_multiplicand[22];
wire w_pp_13_23 = i_multiplier[13] & i_multiplicand[23];
wire w_pp_13_24 = i_multiplier[13] & i_multiplicand[24];
wire w_pp_13_25 = i_multiplier[13] & i_multiplicand[25];
wire w_pp_13_26 = i_multiplier[13] & i_multiplicand[26];
wire w_pp_13_27 = i_multiplier[13] & i_multiplicand[27];
wire w_pp_13_28 = i_multiplier[13] & i_multiplicand[28];
wire w_pp_13_29 = i_multiplier[13] & i_multiplicand[29];
wire w_pp_13_30 = i_multiplier[13] & i_multiplicand[30];
wire w_pp_13_31 = i_multiplier[13] & i_multiplicand[31];
wire w_pp_14_00 = i_multiplier[14] & i_multiplicand[ 0];
wire w_pp_14_01 = i_multiplier[14] & i_multiplicand[ 1];
wire w_pp_14_02 = i_multiplier[14] & i_multiplicand[ 2];
wire w_pp_14_03 = i_multiplier[14] & i_multiplicand[ 3];
wire w_pp_14_04 = i_multiplier[14] & i_multiplicand[ 4];
wire w_pp_14_05 = i_multiplier[14] & i_multiplicand[ 5];
wire w_pp_14_06 = i_multiplier[14] & i_multiplicand[ 6];
wire w_pp_14_07 = i_multiplier[14] & i_multiplicand[ 7];
wire w_pp_14_08 = i_multiplier[14] & i_multiplicand[ 8];
wire w_pp_14_09 = i_multiplier[14] & i_multiplicand[ 9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_14_16 = i_multiplier[14] & i_multiplicand[16];
wire w_pp_14_17 = i_multiplier[14] & i_multiplicand[17];
wire w_pp_14_18 = i_multiplier[14] & i_multiplicand[18];
wire w_pp_14_19 = i_multiplier[14] & i_multiplicand[19];
wire w_pp_14_20 = i_multiplier[14] & i_multiplicand[20];
wire w_pp_14_21 = i_multiplier[14] & i_multiplicand[21];
wire w_pp_14_22 = i_multiplier[14] & i_multiplicand[22];
wire w_pp_14_23 = i_multiplier[14] & i_multiplicand[23];
wire w_pp_14_24 = i_multiplier[14] & i_multiplicand[24];
wire w_pp_14_25 = i_multiplier[14] & i_multiplicand[25];
wire w_pp_14_26 = i_multiplier[14] & i_multiplicand[26];
wire w_pp_14_27 = i_multiplier[14] & i_multiplicand[27];
wire w_pp_14_28 = i_multiplier[14] & i_multiplicand[28];
wire w_pp_14_29 = i_multiplier[14] & i_multiplicand[29];
wire w_pp_14_30 = i_multiplier[14] & i_multiplicand[30];
wire w_pp_14_31 = i_multiplier[14] & i_multiplicand[31];
wire w_pp_15_00 = i_multiplier[15] & i_multiplicand[ 0];
wire w_pp_15_01 = i_multiplier[15] & i_multiplicand[ 1];
wire w_pp_15_02 = i_multiplier[15] & i_multiplicand[ 2];
wire w_pp_15_03 = i_multiplier[15] & i_multiplicand[ 3];
wire w_pp_15_04 = i_multiplier[15] & i_multiplicand[ 4];
wire w_pp_15_05 = i_multiplier[15] & i_multiplicand[ 5];
wire w_pp_15_06 = i_multiplier[15] & i_multiplicand[ 6];
wire w_pp_15_07 = i_multiplier[15] & i_multiplicand[ 7];
wire w_pp_15_08 = i_multiplier[15] & i_multiplicand[ 8];
wire w_pp_15_09 = i_multiplier[15] & i_multiplicand[ 9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];
wire w_pp_15_16 = i_multiplier[15] & i_multiplicand[16];
wire w_pp_15_17 = i_multiplier[15] & i_multiplicand[17];
wire w_pp_15_18 = i_multiplier[15] & i_multiplicand[18];
wire w_pp_15_19 = i_multiplier[15] & i_multiplicand[19];
wire w_pp_15_20 = i_multiplier[15] & i_multiplicand[20];
wire w_pp_15_21 = i_multiplier[15] & i_multiplicand[21];
wire w_pp_15_22 = i_multiplier[15] & i_multiplicand[22];
wire w_pp_15_23 = i_multiplier[15] & i_multiplicand[23];
wire w_pp_15_24 = i_multiplier[15] & i_multiplicand[24];
wire w_pp_15_25 = i_multiplier[15] & i_multiplicand[25];
wire w_pp_15_26 = i_multiplier[15] & i_multiplicand[26];
wire w_pp_15_27 = i_multiplier[15] & i_multiplicand[27];
wire w_pp_15_28 = i_multiplier[15] & i_multiplicand[28];
wire w_pp_15_29 = i_multiplier[15] & i_multiplicand[29];
wire w_pp_15_30 = i_multiplier[15] & i_multiplicand[30];
wire w_pp_15_31 = i_multiplier[15] & i_multiplicand[31];
wire w_pp_16_00 = i_multiplier[16] & i_multiplicand[ 0];
wire w_pp_16_01 = i_multiplier[16] & i_multiplicand[ 1];
wire w_pp_16_02 = i_multiplier[16] & i_multiplicand[ 2];
wire w_pp_16_03 = i_multiplier[16] & i_multiplicand[ 3];
wire w_pp_16_04 = i_multiplier[16] & i_multiplicand[ 4];
wire w_pp_16_05 = i_multiplier[16] & i_multiplicand[ 5];
wire w_pp_16_06 = i_multiplier[16] & i_multiplicand[ 6];
wire w_pp_16_07 = i_multiplier[16] & i_multiplicand[ 7];
wire w_pp_16_08 = i_multiplier[16] & i_multiplicand[ 8];
wire w_pp_16_09 = i_multiplier[16] & i_multiplicand[ 9];
wire w_pp_16_10 = i_multiplier[16] & i_multiplicand[10];
wire w_pp_16_11 = i_multiplier[16] & i_multiplicand[11];
wire w_pp_16_12 = i_multiplier[16] & i_multiplicand[12];
wire w_pp_16_13 = i_multiplier[16] & i_multiplicand[13];
wire w_pp_16_14 = i_multiplier[16] & i_multiplicand[14];
wire w_pp_16_15 = i_multiplier[16] & i_multiplicand[15];
wire w_pp_16_16 = i_multiplier[16] & i_multiplicand[16];
wire w_pp_16_17 = i_multiplier[16] & i_multiplicand[17];
wire w_pp_16_18 = i_multiplier[16] & i_multiplicand[18];
wire w_pp_16_19 = i_multiplier[16] & i_multiplicand[19];
wire w_pp_16_20 = i_multiplier[16] & i_multiplicand[20];
wire w_pp_16_21 = i_multiplier[16] & i_multiplicand[21];
wire w_pp_16_22 = i_multiplier[16] & i_multiplicand[22];
wire w_pp_16_23 = i_multiplier[16] & i_multiplicand[23];
wire w_pp_16_24 = i_multiplier[16] & i_multiplicand[24];
wire w_pp_16_25 = i_multiplier[16] & i_multiplicand[25];
wire w_pp_16_26 = i_multiplier[16] & i_multiplicand[26];
wire w_pp_16_27 = i_multiplier[16] & i_multiplicand[27];
wire w_pp_16_28 = i_multiplier[16] & i_multiplicand[28];
wire w_pp_16_29 = i_multiplier[16] & i_multiplicand[29];
wire w_pp_16_30 = i_multiplier[16] & i_multiplicand[30];
wire w_pp_16_31 = i_multiplier[16] & i_multiplicand[31];
wire w_pp_17_00 = i_multiplier[17] & i_multiplicand[ 0];
wire w_pp_17_01 = i_multiplier[17] & i_multiplicand[ 1];
wire w_pp_17_02 = i_multiplier[17] & i_multiplicand[ 2];
wire w_pp_17_03 = i_multiplier[17] & i_multiplicand[ 3];
wire w_pp_17_04 = i_multiplier[17] & i_multiplicand[ 4];
wire w_pp_17_05 = i_multiplier[17] & i_multiplicand[ 5];
wire w_pp_17_06 = i_multiplier[17] & i_multiplicand[ 6];
wire w_pp_17_07 = i_multiplier[17] & i_multiplicand[ 7];
wire w_pp_17_08 = i_multiplier[17] & i_multiplicand[ 8];
wire w_pp_17_09 = i_multiplier[17] & i_multiplicand[ 9];
wire w_pp_17_10 = i_multiplier[17] & i_multiplicand[10];
wire w_pp_17_11 = i_multiplier[17] & i_multiplicand[11];
wire w_pp_17_12 = i_multiplier[17] & i_multiplicand[12];
wire w_pp_17_13 = i_multiplier[17] & i_multiplicand[13];
wire w_pp_17_14 = i_multiplier[17] & i_multiplicand[14];
wire w_pp_17_15 = i_multiplier[17] & i_multiplicand[15];
wire w_pp_17_16 = i_multiplier[17] & i_multiplicand[16];
wire w_pp_17_17 = i_multiplier[17] & i_multiplicand[17];
wire w_pp_17_18 = i_multiplier[17] & i_multiplicand[18];
wire w_pp_17_19 = i_multiplier[17] & i_multiplicand[19];
wire w_pp_17_20 = i_multiplier[17] & i_multiplicand[20];
wire w_pp_17_21 = i_multiplier[17] & i_multiplicand[21];
wire w_pp_17_22 = i_multiplier[17] & i_multiplicand[22];
wire w_pp_17_23 = i_multiplier[17] & i_multiplicand[23];
wire w_pp_17_24 = i_multiplier[17] & i_multiplicand[24];
wire w_pp_17_25 = i_multiplier[17] & i_multiplicand[25];
wire w_pp_17_26 = i_multiplier[17] & i_multiplicand[26];
wire w_pp_17_27 = i_multiplier[17] & i_multiplicand[27];
wire w_pp_17_28 = i_multiplier[17] & i_multiplicand[28];
wire w_pp_17_29 = i_multiplier[17] & i_multiplicand[29];
wire w_pp_17_30 = i_multiplier[17] & i_multiplicand[30];
wire w_pp_17_31 = i_multiplier[17] & i_multiplicand[31];
wire w_pp_18_00 = i_multiplier[18] & i_multiplicand[ 0];
wire w_pp_18_01 = i_multiplier[18] & i_multiplicand[ 1];
wire w_pp_18_02 = i_multiplier[18] & i_multiplicand[ 2];
wire w_pp_18_03 = i_multiplier[18] & i_multiplicand[ 3];
wire w_pp_18_04 = i_multiplier[18] & i_multiplicand[ 4];
wire w_pp_18_05 = i_multiplier[18] & i_multiplicand[ 5];
wire w_pp_18_06 = i_multiplier[18] & i_multiplicand[ 6];
wire w_pp_18_07 = i_multiplier[18] & i_multiplicand[ 7];
wire w_pp_18_08 = i_multiplier[18] & i_multiplicand[ 8];
wire w_pp_18_09 = i_multiplier[18] & i_multiplicand[ 9];
wire w_pp_18_10 = i_multiplier[18] & i_multiplicand[10];
wire w_pp_18_11 = i_multiplier[18] & i_multiplicand[11];
wire w_pp_18_12 = i_multiplier[18] & i_multiplicand[12];
wire w_pp_18_13 = i_multiplier[18] & i_multiplicand[13];
wire w_pp_18_14 = i_multiplier[18] & i_multiplicand[14];
wire w_pp_18_15 = i_multiplier[18] & i_multiplicand[15];
wire w_pp_18_16 = i_multiplier[18] & i_multiplicand[16];
wire w_pp_18_17 = i_multiplier[18] & i_multiplicand[17];
wire w_pp_18_18 = i_multiplier[18] & i_multiplicand[18];
wire w_pp_18_19 = i_multiplier[18] & i_multiplicand[19];
wire w_pp_18_20 = i_multiplier[18] & i_multiplicand[20];
wire w_pp_18_21 = i_multiplier[18] & i_multiplicand[21];
wire w_pp_18_22 = i_multiplier[18] & i_multiplicand[22];
wire w_pp_18_23 = i_multiplier[18] & i_multiplicand[23];
wire w_pp_18_24 = i_multiplier[18] & i_multiplicand[24];
wire w_pp_18_25 = i_multiplier[18] & i_multiplicand[25];
wire w_pp_18_26 = i_multiplier[18] & i_multiplicand[26];
wire w_pp_18_27 = i_multiplier[18] & i_multiplicand[27];
wire w_pp_18_28 = i_multiplier[18] & i_multiplicand[28];
wire w_pp_18_29 = i_multiplier[18] & i_multiplicand[29];
wire w_pp_18_30 = i_multiplier[18] & i_multiplicand[30];
wire w_pp_18_31 = i_multiplier[18] & i_multiplicand[31];
wire w_pp_19_00 = i_multiplier[19] & i_multiplicand[ 0];
wire w_pp_19_01 = i_multiplier[19] & i_multiplicand[ 1];
wire w_pp_19_02 = i_multiplier[19] & i_multiplicand[ 2];
wire w_pp_19_03 = i_multiplier[19] & i_multiplicand[ 3];
wire w_pp_19_04 = i_multiplier[19] & i_multiplicand[ 4];
wire w_pp_19_05 = i_multiplier[19] & i_multiplicand[ 5];
wire w_pp_19_06 = i_multiplier[19] & i_multiplicand[ 6];
wire w_pp_19_07 = i_multiplier[19] & i_multiplicand[ 7];
wire w_pp_19_08 = i_multiplier[19] & i_multiplicand[ 8];
wire w_pp_19_09 = i_multiplier[19] & i_multiplicand[ 9];
wire w_pp_19_10 = i_multiplier[19] & i_multiplicand[10];
wire w_pp_19_11 = i_multiplier[19] & i_multiplicand[11];
wire w_pp_19_12 = i_multiplier[19] & i_multiplicand[12];
wire w_pp_19_13 = i_multiplier[19] & i_multiplicand[13];
wire w_pp_19_14 = i_multiplier[19] & i_multiplicand[14];
wire w_pp_19_15 = i_multiplier[19] & i_multiplicand[15];
wire w_pp_19_16 = i_multiplier[19] & i_multiplicand[16];
wire w_pp_19_17 = i_multiplier[19] & i_multiplicand[17];
wire w_pp_19_18 = i_multiplier[19] & i_multiplicand[18];
wire w_pp_19_19 = i_multiplier[19] & i_multiplicand[19];
wire w_pp_19_20 = i_multiplier[19] & i_multiplicand[20];
wire w_pp_19_21 = i_multiplier[19] & i_multiplicand[21];
wire w_pp_19_22 = i_multiplier[19] & i_multiplicand[22];
wire w_pp_19_23 = i_multiplier[19] & i_multiplicand[23];
wire w_pp_19_24 = i_multiplier[19] & i_multiplicand[24];
wire w_pp_19_25 = i_multiplier[19] & i_multiplicand[25];
wire w_pp_19_26 = i_multiplier[19] & i_multiplicand[26];
wire w_pp_19_27 = i_multiplier[19] & i_multiplicand[27];
wire w_pp_19_28 = i_multiplier[19] & i_multiplicand[28];
wire w_pp_19_29 = i_multiplier[19] & i_multiplicand[29];
wire w_pp_19_30 = i_multiplier[19] & i_multiplicand[30];
wire w_pp_19_31 = i_multiplier[19] & i_multiplicand[31];
wire w_pp_20_00 = i_multiplier[20] & i_multiplicand[ 0];
wire w_pp_20_01 = i_multiplier[20] & i_multiplicand[ 1];
wire w_pp_20_02 = i_multiplier[20] & i_multiplicand[ 2];
wire w_pp_20_03 = i_multiplier[20] & i_multiplicand[ 3];
wire w_pp_20_04 = i_multiplier[20] & i_multiplicand[ 4];
wire w_pp_20_05 = i_multiplier[20] & i_multiplicand[ 5];
wire w_pp_20_06 = i_multiplier[20] & i_multiplicand[ 6];
wire w_pp_20_07 = i_multiplier[20] & i_multiplicand[ 7];
wire w_pp_20_08 = i_multiplier[20] & i_multiplicand[ 8];
wire w_pp_20_09 = i_multiplier[20] & i_multiplicand[ 9];
wire w_pp_20_10 = i_multiplier[20] & i_multiplicand[10];
wire w_pp_20_11 = i_multiplier[20] & i_multiplicand[11];
wire w_pp_20_12 = i_multiplier[20] & i_multiplicand[12];
wire w_pp_20_13 = i_multiplier[20] & i_multiplicand[13];
wire w_pp_20_14 = i_multiplier[20] & i_multiplicand[14];
wire w_pp_20_15 = i_multiplier[20] & i_multiplicand[15];
wire w_pp_20_16 = i_multiplier[20] & i_multiplicand[16];
wire w_pp_20_17 = i_multiplier[20] & i_multiplicand[17];
wire w_pp_20_18 = i_multiplier[20] & i_multiplicand[18];
wire w_pp_20_19 = i_multiplier[20] & i_multiplicand[19];
wire w_pp_20_20 = i_multiplier[20] & i_multiplicand[20];
wire w_pp_20_21 = i_multiplier[20] & i_multiplicand[21];
wire w_pp_20_22 = i_multiplier[20] & i_multiplicand[22];
wire w_pp_20_23 = i_multiplier[20] & i_multiplicand[23];
wire w_pp_20_24 = i_multiplier[20] & i_multiplicand[24];
wire w_pp_20_25 = i_multiplier[20] & i_multiplicand[25];
wire w_pp_20_26 = i_multiplier[20] & i_multiplicand[26];
wire w_pp_20_27 = i_multiplier[20] & i_multiplicand[27];
wire w_pp_20_28 = i_multiplier[20] & i_multiplicand[28];
wire w_pp_20_29 = i_multiplier[20] & i_multiplicand[29];
wire w_pp_20_30 = i_multiplier[20] & i_multiplicand[30];
wire w_pp_20_31 = i_multiplier[20] & i_multiplicand[31];
wire w_pp_21_00 = i_multiplier[21] & i_multiplicand[ 0];
wire w_pp_21_01 = i_multiplier[21] & i_multiplicand[ 1];
wire w_pp_21_02 = i_multiplier[21] & i_multiplicand[ 2];
wire w_pp_21_03 = i_multiplier[21] & i_multiplicand[ 3];
wire w_pp_21_04 = i_multiplier[21] & i_multiplicand[ 4];
wire w_pp_21_05 = i_multiplier[21] & i_multiplicand[ 5];
wire w_pp_21_06 = i_multiplier[21] & i_multiplicand[ 6];
wire w_pp_21_07 = i_multiplier[21] & i_multiplicand[ 7];
wire w_pp_21_08 = i_multiplier[21] & i_multiplicand[ 8];
wire w_pp_21_09 = i_multiplier[21] & i_multiplicand[ 9];
wire w_pp_21_10 = i_multiplier[21] & i_multiplicand[10];
wire w_pp_21_11 = i_multiplier[21] & i_multiplicand[11];
wire w_pp_21_12 = i_multiplier[21] & i_multiplicand[12];
wire w_pp_21_13 = i_multiplier[21] & i_multiplicand[13];
wire w_pp_21_14 = i_multiplier[21] & i_multiplicand[14];
wire w_pp_21_15 = i_multiplier[21] & i_multiplicand[15];
wire w_pp_21_16 = i_multiplier[21] & i_multiplicand[16];
wire w_pp_21_17 = i_multiplier[21] & i_multiplicand[17];
wire w_pp_21_18 = i_multiplier[21] & i_multiplicand[18];
wire w_pp_21_19 = i_multiplier[21] & i_multiplicand[19];
wire w_pp_21_20 = i_multiplier[21] & i_multiplicand[20];
wire w_pp_21_21 = i_multiplier[21] & i_multiplicand[21];
wire w_pp_21_22 = i_multiplier[21] & i_multiplicand[22];
wire w_pp_21_23 = i_multiplier[21] & i_multiplicand[23];
wire w_pp_21_24 = i_multiplier[21] & i_multiplicand[24];
wire w_pp_21_25 = i_multiplier[21] & i_multiplicand[25];
wire w_pp_21_26 = i_multiplier[21] & i_multiplicand[26];
wire w_pp_21_27 = i_multiplier[21] & i_multiplicand[27];
wire w_pp_21_28 = i_multiplier[21] & i_multiplicand[28];
wire w_pp_21_29 = i_multiplier[21] & i_multiplicand[29];
wire w_pp_21_30 = i_multiplier[21] & i_multiplicand[30];
wire w_pp_21_31 = i_multiplier[21] & i_multiplicand[31];
wire w_pp_22_00 = i_multiplier[22] & i_multiplicand[ 0];
wire w_pp_22_01 = i_multiplier[22] & i_multiplicand[ 1];
wire w_pp_22_02 = i_multiplier[22] & i_multiplicand[ 2];
wire w_pp_22_03 = i_multiplier[22] & i_multiplicand[ 3];
wire w_pp_22_04 = i_multiplier[22] & i_multiplicand[ 4];
wire w_pp_22_05 = i_multiplier[22] & i_multiplicand[ 5];
wire w_pp_22_06 = i_multiplier[22] & i_multiplicand[ 6];
wire w_pp_22_07 = i_multiplier[22] & i_multiplicand[ 7];
wire w_pp_22_08 = i_multiplier[22] & i_multiplicand[ 8];
wire w_pp_22_09 = i_multiplier[22] & i_multiplicand[ 9];
wire w_pp_22_10 = i_multiplier[22] & i_multiplicand[10];
wire w_pp_22_11 = i_multiplier[22] & i_multiplicand[11];
wire w_pp_22_12 = i_multiplier[22] & i_multiplicand[12];
wire w_pp_22_13 = i_multiplier[22] & i_multiplicand[13];
wire w_pp_22_14 = i_multiplier[22] & i_multiplicand[14];
wire w_pp_22_15 = i_multiplier[22] & i_multiplicand[15];
wire w_pp_22_16 = i_multiplier[22] & i_multiplicand[16];
wire w_pp_22_17 = i_multiplier[22] & i_multiplicand[17];
wire w_pp_22_18 = i_multiplier[22] & i_multiplicand[18];
wire w_pp_22_19 = i_multiplier[22] & i_multiplicand[19];
wire w_pp_22_20 = i_multiplier[22] & i_multiplicand[20];
wire w_pp_22_21 = i_multiplier[22] & i_multiplicand[21];
wire w_pp_22_22 = i_multiplier[22] & i_multiplicand[22];
wire w_pp_22_23 = i_multiplier[22] & i_multiplicand[23];
wire w_pp_22_24 = i_multiplier[22] & i_multiplicand[24];
wire w_pp_22_25 = i_multiplier[22] & i_multiplicand[25];
wire w_pp_22_26 = i_multiplier[22] & i_multiplicand[26];
wire w_pp_22_27 = i_multiplier[22] & i_multiplicand[27];
wire w_pp_22_28 = i_multiplier[22] & i_multiplicand[28];
wire w_pp_22_29 = i_multiplier[22] & i_multiplicand[29];
wire w_pp_22_30 = i_multiplier[22] & i_multiplicand[30];
wire w_pp_22_31 = i_multiplier[22] & i_multiplicand[31];
wire w_pp_23_00 = i_multiplier[23] & i_multiplicand[ 0];
wire w_pp_23_01 = i_multiplier[23] & i_multiplicand[ 1];
wire w_pp_23_02 = i_multiplier[23] & i_multiplicand[ 2];
wire w_pp_23_03 = i_multiplier[23] & i_multiplicand[ 3];
wire w_pp_23_04 = i_multiplier[23] & i_multiplicand[ 4];
wire w_pp_23_05 = i_multiplier[23] & i_multiplicand[ 5];
wire w_pp_23_06 = i_multiplier[23] & i_multiplicand[ 6];
wire w_pp_23_07 = i_multiplier[23] & i_multiplicand[ 7];
wire w_pp_23_08 = i_multiplier[23] & i_multiplicand[ 8];
wire w_pp_23_09 = i_multiplier[23] & i_multiplicand[ 9];
wire w_pp_23_10 = i_multiplier[23] & i_multiplicand[10];
wire w_pp_23_11 = i_multiplier[23] & i_multiplicand[11];
wire w_pp_23_12 = i_multiplier[23] & i_multiplicand[12];
wire w_pp_23_13 = i_multiplier[23] & i_multiplicand[13];
wire w_pp_23_14 = i_multiplier[23] & i_multiplicand[14];
wire w_pp_23_15 = i_multiplier[23] & i_multiplicand[15];
wire w_pp_23_16 = i_multiplier[23] & i_multiplicand[16];
wire w_pp_23_17 = i_multiplier[23] & i_multiplicand[17];
wire w_pp_23_18 = i_multiplier[23] & i_multiplicand[18];
wire w_pp_23_19 = i_multiplier[23] & i_multiplicand[19];
wire w_pp_23_20 = i_multiplier[23] & i_multiplicand[20];
wire w_pp_23_21 = i_multiplier[23] & i_multiplicand[21];
wire w_pp_23_22 = i_multiplier[23] & i_multiplicand[22];
wire w_pp_23_23 = i_multiplier[23] & i_multiplicand[23];
wire w_pp_23_24 = i_multiplier[23] & i_multiplicand[24];
wire w_pp_23_25 = i_multiplier[23] & i_multiplicand[25];
wire w_pp_23_26 = i_multiplier[23] & i_multiplicand[26];
wire w_pp_23_27 = i_multiplier[23] & i_multiplicand[27];
wire w_pp_23_28 = i_multiplier[23] & i_multiplicand[28];
wire w_pp_23_29 = i_multiplier[23] & i_multiplicand[29];
wire w_pp_23_30 = i_multiplier[23] & i_multiplicand[30];
wire w_pp_23_31 = i_multiplier[23] & i_multiplicand[31];
wire w_pp_24_00 = i_multiplier[24] & i_multiplicand[ 0];
wire w_pp_24_01 = i_multiplier[24] & i_multiplicand[ 1];
wire w_pp_24_02 = i_multiplier[24] & i_multiplicand[ 2];
wire w_pp_24_03 = i_multiplier[24] & i_multiplicand[ 3];
wire w_pp_24_04 = i_multiplier[24] & i_multiplicand[ 4];
wire w_pp_24_05 = i_multiplier[24] & i_multiplicand[ 5];
wire w_pp_24_06 = i_multiplier[24] & i_multiplicand[ 6];
wire w_pp_24_07 = i_multiplier[24] & i_multiplicand[ 7];
wire w_pp_24_08 = i_multiplier[24] & i_multiplicand[ 8];
wire w_pp_24_09 = i_multiplier[24] & i_multiplicand[ 9];
wire w_pp_24_10 = i_multiplier[24] & i_multiplicand[10];
wire w_pp_24_11 = i_multiplier[24] & i_multiplicand[11];
wire w_pp_24_12 = i_multiplier[24] & i_multiplicand[12];
wire w_pp_24_13 = i_multiplier[24] & i_multiplicand[13];
wire w_pp_24_14 = i_multiplier[24] & i_multiplicand[14];
wire w_pp_24_15 = i_multiplier[24] & i_multiplicand[15];
wire w_pp_24_16 = i_multiplier[24] & i_multiplicand[16];
wire w_pp_24_17 = i_multiplier[24] & i_multiplicand[17];
wire w_pp_24_18 = i_multiplier[24] & i_multiplicand[18];
wire w_pp_24_19 = i_multiplier[24] & i_multiplicand[19];
wire w_pp_24_20 = i_multiplier[24] & i_multiplicand[20];
wire w_pp_24_21 = i_multiplier[24] & i_multiplicand[21];
wire w_pp_24_22 = i_multiplier[24] & i_multiplicand[22];
wire w_pp_24_23 = i_multiplier[24] & i_multiplicand[23];
wire w_pp_24_24 = i_multiplier[24] & i_multiplicand[24];
wire w_pp_24_25 = i_multiplier[24] & i_multiplicand[25];
wire w_pp_24_26 = i_multiplier[24] & i_multiplicand[26];
wire w_pp_24_27 = i_multiplier[24] & i_multiplicand[27];
wire w_pp_24_28 = i_multiplier[24] & i_multiplicand[28];
wire w_pp_24_29 = i_multiplier[24] & i_multiplicand[29];
wire w_pp_24_30 = i_multiplier[24] & i_multiplicand[30];
wire w_pp_24_31 = i_multiplier[24] & i_multiplicand[31];
wire w_pp_25_00 = i_multiplier[25] & i_multiplicand[ 0];
wire w_pp_25_01 = i_multiplier[25] & i_multiplicand[ 1];
wire w_pp_25_02 = i_multiplier[25] & i_multiplicand[ 2];
wire w_pp_25_03 = i_multiplier[25] & i_multiplicand[ 3];
wire w_pp_25_04 = i_multiplier[25] & i_multiplicand[ 4];
wire w_pp_25_05 = i_multiplier[25] & i_multiplicand[ 5];
wire w_pp_25_06 = i_multiplier[25] & i_multiplicand[ 6];
wire w_pp_25_07 = i_multiplier[25] & i_multiplicand[ 7];
wire w_pp_25_08 = i_multiplier[25] & i_multiplicand[ 8];
wire w_pp_25_09 = i_multiplier[25] & i_multiplicand[ 9];
wire w_pp_25_10 = i_multiplier[25] & i_multiplicand[10];
wire w_pp_25_11 = i_multiplier[25] & i_multiplicand[11];
wire w_pp_25_12 = i_multiplier[25] & i_multiplicand[12];
wire w_pp_25_13 = i_multiplier[25] & i_multiplicand[13];
wire w_pp_25_14 = i_multiplier[25] & i_multiplicand[14];
wire w_pp_25_15 = i_multiplier[25] & i_multiplicand[15];
wire w_pp_25_16 = i_multiplier[25] & i_multiplicand[16];
wire w_pp_25_17 = i_multiplier[25] & i_multiplicand[17];
wire w_pp_25_18 = i_multiplier[25] & i_multiplicand[18];
wire w_pp_25_19 = i_multiplier[25] & i_multiplicand[19];
wire w_pp_25_20 = i_multiplier[25] & i_multiplicand[20];
wire w_pp_25_21 = i_multiplier[25] & i_multiplicand[21];
wire w_pp_25_22 = i_multiplier[25] & i_multiplicand[22];
wire w_pp_25_23 = i_multiplier[25] & i_multiplicand[23];
wire w_pp_25_24 = i_multiplier[25] & i_multiplicand[24];
wire w_pp_25_25 = i_multiplier[25] & i_multiplicand[25];
wire w_pp_25_26 = i_multiplier[25] & i_multiplicand[26];
wire w_pp_25_27 = i_multiplier[25] & i_multiplicand[27];
wire w_pp_25_28 = i_multiplier[25] & i_multiplicand[28];
wire w_pp_25_29 = i_multiplier[25] & i_multiplicand[29];
wire w_pp_25_30 = i_multiplier[25] & i_multiplicand[30];
wire w_pp_25_31 = i_multiplier[25] & i_multiplicand[31];
wire w_pp_26_00 = i_multiplier[26] & i_multiplicand[ 0];
wire w_pp_26_01 = i_multiplier[26] & i_multiplicand[ 1];
wire w_pp_26_02 = i_multiplier[26] & i_multiplicand[ 2];
wire w_pp_26_03 = i_multiplier[26] & i_multiplicand[ 3];
wire w_pp_26_04 = i_multiplier[26] & i_multiplicand[ 4];
wire w_pp_26_05 = i_multiplier[26] & i_multiplicand[ 5];
wire w_pp_26_06 = i_multiplier[26] & i_multiplicand[ 6];
wire w_pp_26_07 = i_multiplier[26] & i_multiplicand[ 7];
wire w_pp_26_08 = i_multiplier[26] & i_multiplicand[ 8];
wire w_pp_26_09 = i_multiplier[26] & i_multiplicand[ 9];
wire w_pp_26_10 = i_multiplier[26] & i_multiplicand[10];
wire w_pp_26_11 = i_multiplier[26] & i_multiplicand[11];
wire w_pp_26_12 = i_multiplier[26] & i_multiplicand[12];
wire w_pp_26_13 = i_multiplier[26] & i_multiplicand[13];
wire w_pp_26_14 = i_multiplier[26] & i_multiplicand[14];
wire w_pp_26_15 = i_multiplier[26] & i_multiplicand[15];
wire w_pp_26_16 = i_multiplier[26] & i_multiplicand[16];
wire w_pp_26_17 = i_multiplier[26] & i_multiplicand[17];
wire w_pp_26_18 = i_multiplier[26] & i_multiplicand[18];
wire w_pp_26_19 = i_multiplier[26] & i_multiplicand[19];
wire w_pp_26_20 = i_multiplier[26] & i_multiplicand[20];
wire w_pp_26_21 = i_multiplier[26] & i_multiplicand[21];
wire w_pp_26_22 = i_multiplier[26] & i_multiplicand[22];
wire w_pp_26_23 = i_multiplier[26] & i_multiplicand[23];
wire w_pp_26_24 = i_multiplier[26] & i_multiplicand[24];
wire w_pp_26_25 = i_multiplier[26] & i_multiplicand[25];
wire w_pp_26_26 = i_multiplier[26] & i_multiplicand[26];
wire w_pp_26_27 = i_multiplier[26] & i_multiplicand[27];
wire w_pp_26_28 = i_multiplier[26] & i_multiplicand[28];
wire w_pp_26_29 = i_multiplier[26] & i_multiplicand[29];
wire w_pp_26_30 = i_multiplier[26] & i_multiplicand[30];
wire w_pp_26_31 = i_multiplier[26] & i_multiplicand[31];
wire w_pp_27_00 = i_multiplier[27] & i_multiplicand[ 0];
wire w_pp_27_01 = i_multiplier[27] & i_multiplicand[ 1];
wire w_pp_27_02 = i_multiplier[27] & i_multiplicand[ 2];
wire w_pp_27_03 = i_multiplier[27] & i_multiplicand[ 3];
wire w_pp_27_04 = i_multiplier[27] & i_multiplicand[ 4];
wire w_pp_27_05 = i_multiplier[27] & i_multiplicand[ 5];
wire w_pp_27_06 = i_multiplier[27] & i_multiplicand[ 6];
wire w_pp_27_07 = i_multiplier[27] & i_multiplicand[ 7];
wire w_pp_27_08 = i_multiplier[27] & i_multiplicand[ 8];
wire w_pp_27_09 = i_multiplier[27] & i_multiplicand[ 9];
wire w_pp_27_10 = i_multiplier[27] & i_multiplicand[10];
wire w_pp_27_11 = i_multiplier[27] & i_multiplicand[11];
wire w_pp_27_12 = i_multiplier[27] & i_multiplicand[12];
wire w_pp_27_13 = i_multiplier[27] & i_multiplicand[13];
wire w_pp_27_14 = i_multiplier[27] & i_multiplicand[14];
wire w_pp_27_15 = i_multiplier[27] & i_multiplicand[15];
wire w_pp_27_16 = i_multiplier[27] & i_multiplicand[16];
wire w_pp_27_17 = i_multiplier[27] & i_multiplicand[17];
wire w_pp_27_18 = i_multiplier[27] & i_multiplicand[18];
wire w_pp_27_19 = i_multiplier[27] & i_multiplicand[19];
wire w_pp_27_20 = i_multiplier[27] & i_multiplicand[20];
wire w_pp_27_21 = i_multiplier[27] & i_multiplicand[21];
wire w_pp_27_22 = i_multiplier[27] & i_multiplicand[22];
wire w_pp_27_23 = i_multiplier[27] & i_multiplicand[23];
wire w_pp_27_24 = i_multiplier[27] & i_multiplicand[24];
wire w_pp_27_25 = i_multiplier[27] & i_multiplicand[25];
wire w_pp_27_26 = i_multiplier[27] & i_multiplicand[26];
wire w_pp_27_27 = i_multiplier[27] & i_multiplicand[27];
wire w_pp_27_28 = i_multiplier[27] & i_multiplicand[28];
wire w_pp_27_29 = i_multiplier[27] & i_multiplicand[29];
wire w_pp_27_30 = i_multiplier[27] & i_multiplicand[30];
wire w_pp_27_31 = i_multiplier[27] & i_multiplicand[31];
wire w_pp_28_00 = i_multiplier[28] & i_multiplicand[ 0];
wire w_pp_28_01 = i_multiplier[28] & i_multiplicand[ 1];
wire w_pp_28_02 = i_multiplier[28] & i_multiplicand[ 2];
wire w_pp_28_03 = i_multiplier[28] & i_multiplicand[ 3];
wire w_pp_28_04 = i_multiplier[28] & i_multiplicand[ 4];
wire w_pp_28_05 = i_multiplier[28] & i_multiplicand[ 5];
wire w_pp_28_06 = i_multiplier[28] & i_multiplicand[ 6];
wire w_pp_28_07 = i_multiplier[28] & i_multiplicand[ 7];
wire w_pp_28_08 = i_multiplier[28] & i_multiplicand[ 8];
wire w_pp_28_09 = i_multiplier[28] & i_multiplicand[ 9];
wire w_pp_28_10 = i_multiplier[28] & i_multiplicand[10];
wire w_pp_28_11 = i_multiplier[28] & i_multiplicand[11];
wire w_pp_28_12 = i_multiplier[28] & i_multiplicand[12];
wire w_pp_28_13 = i_multiplier[28] & i_multiplicand[13];
wire w_pp_28_14 = i_multiplier[28] & i_multiplicand[14];
wire w_pp_28_15 = i_multiplier[28] & i_multiplicand[15];
wire w_pp_28_16 = i_multiplier[28] & i_multiplicand[16];
wire w_pp_28_17 = i_multiplier[28] & i_multiplicand[17];
wire w_pp_28_18 = i_multiplier[28] & i_multiplicand[18];
wire w_pp_28_19 = i_multiplier[28] & i_multiplicand[19];
wire w_pp_28_20 = i_multiplier[28] & i_multiplicand[20];
wire w_pp_28_21 = i_multiplier[28] & i_multiplicand[21];
wire w_pp_28_22 = i_multiplier[28] & i_multiplicand[22];
wire w_pp_28_23 = i_multiplier[28] & i_multiplicand[23];
wire w_pp_28_24 = i_multiplier[28] & i_multiplicand[24];
wire w_pp_28_25 = i_multiplier[28] & i_multiplicand[25];
wire w_pp_28_26 = i_multiplier[28] & i_multiplicand[26];
wire w_pp_28_27 = i_multiplier[28] & i_multiplicand[27];
wire w_pp_28_28 = i_multiplier[28] & i_multiplicand[28];
wire w_pp_28_29 = i_multiplier[28] & i_multiplicand[29];
wire w_pp_28_30 = i_multiplier[28] & i_multiplicand[30];
wire w_pp_28_31 = i_multiplier[28] & i_multiplicand[31];
wire w_pp_29_00 = i_multiplier[29] & i_multiplicand[ 0];
wire w_pp_29_01 = i_multiplier[29] & i_multiplicand[ 1];
wire w_pp_29_02 = i_multiplier[29] & i_multiplicand[ 2];
wire w_pp_29_03 = i_multiplier[29] & i_multiplicand[ 3];
wire w_pp_29_04 = i_multiplier[29] & i_multiplicand[ 4];
wire w_pp_29_05 = i_multiplier[29] & i_multiplicand[ 5];
wire w_pp_29_06 = i_multiplier[29] & i_multiplicand[ 6];
wire w_pp_29_07 = i_multiplier[29] & i_multiplicand[ 7];
wire w_pp_29_08 = i_multiplier[29] & i_multiplicand[ 8];
wire w_pp_29_09 = i_multiplier[29] & i_multiplicand[ 9];
wire w_pp_29_10 = i_multiplier[29] & i_multiplicand[10];
wire w_pp_29_11 = i_multiplier[29] & i_multiplicand[11];
wire w_pp_29_12 = i_multiplier[29] & i_multiplicand[12];
wire w_pp_29_13 = i_multiplier[29] & i_multiplicand[13];
wire w_pp_29_14 = i_multiplier[29] & i_multiplicand[14];
wire w_pp_29_15 = i_multiplier[29] & i_multiplicand[15];
wire w_pp_29_16 = i_multiplier[29] & i_multiplicand[16];
wire w_pp_29_17 = i_multiplier[29] & i_multiplicand[17];
wire w_pp_29_18 = i_multiplier[29] & i_multiplicand[18];
wire w_pp_29_19 = i_multiplier[29] & i_multiplicand[19];
wire w_pp_29_20 = i_multiplier[29] & i_multiplicand[20];
wire w_pp_29_21 = i_multiplier[29] & i_multiplicand[21];
wire w_pp_29_22 = i_multiplier[29] & i_multiplicand[22];
wire w_pp_29_23 = i_multiplier[29] & i_multiplicand[23];
wire w_pp_29_24 = i_multiplier[29] & i_multiplicand[24];
wire w_pp_29_25 = i_multiplier[29] & i_multiplicand[25];
wire w_pp_29_26 = i_multiplier[29] & i_multiplicand[26];
wire w_pp_29_27 = i_multiplier[29] & i_multiplicand[27];
wire w_pp_29_28 = i_multiplier[29] & i_multiplicand[28];
wire w_pp_29_29 = i_multiplier[29] & i_multiplicand[29];
wire w_pp_29_30 = i_multiplier[29] & i_multiplicand[30];
wire w_pp_29_31 = i_multiplier[29] & i_multiplicand[31];
wire w_pp_30_00 = i_multiplier[30] & i_multiplicand[ 0];
wire w_pp_30_01 = i_multiplier[30] & i_multiplicand[ 1];
wire w_pp_30_02 = i_multiplier[30] & i_multiplicand[ 2];
wire w_pp_30_03 = i_multiplier[30] & i_multiplicand[ 3];
wire w_pp_30_04 = i_multiplier[30] & i_multiplicand[ 4];
wire w_pp_30_05 = i_multiplier[30] & i_multiplicand[ 5];
wire w_pp_30_06 = i_multiplier[30] & i_multiplicand[ 6];
wire w_pp_30_07 = i_multiplier[30] & i_multiplicand[ 7];
wire w_pp_30_08 = i_multiplier[30] & i_multiplicand[ 8];
wire w_pp_30_09 = i_multiplier[30] & i_multiplicand[ 9];
wire w_pp_30_10 = i_multiplier[30] & i_multiplicand[10];
wire w_pp_30_11 = i_multiplier[30] & i_multiplicand[11];
wire w_pp_30_12 = i_multiplier[30] & i_multiplicand[12];
wire w_pp_30_13 = i_multiplier[30] & i_multiplicand[13];
wire w_pp_30_14 = i_multiplier[30] & i_multiplicand[14];
wire w_pp_30_15 = i_multiplier[30] & i_multiplicand[15];
wire w_pp_30_16 = i_multiplier[30] & i_multiplicand[16];
wire w_pp_30_17 = i_multiplier[30] & i_multiplicand[17];
wire w_pp_30_18 = i_multiplier[30] & i_multiplicand[18];
wire w_pp_30_19 = i_multiplier[30] & i_multiplicand[19];
wire w_pp_30_20 = i_multiplier[30] & i_multiplicand[20];
wire w_pp_30_21 = i_multiplier[30] & i_multiplicand[21];
wire w_pp_30_22 = i_multiplier[30] & i_multiplicand[22];
wire w_pp_30_23 = i_multiplier[30] & i_multiplicand[23];
wire w_pp_30_24 = i_multiplier[30] & i_multiplicand[24];
wire w_pp_30_25 = i_multiplier[30] & i_multiplicand[25];
wire w_pp_30_26 = i_multiplier[30] & i_multiplicand[26];
wire w_pp_30_27 = i_multiplier[30] & i_multiplicand[27];
wire w_pp_30_28 = i_multiplier[30] & i_multiplicand[28];
wire w_pp_30_29 = i_multiplier[30] & i_multiplicand[29];
wire w_pp_30_30 = i_multiplier[30] & i_multiplicand[30];
wire w_pp_30_31 = i_multiplier[30] & i_multiplicand[31];
wire w_pp_31_00 = i_multiplier[31] & i_multiplicand[ 0];
wire w_pp_31_01 = i_multiplier[31] & i_multiplicand[ 1];
wire w_pp_31_02 = i_multiplier[31] & i_multiplicand[ 2];
wire w_pp_31_03 = i_multiplier[31] & i_multiplicand[ 3];
wire w_pp_31_04 = i_multiplier[31] & i_multiplicand[ 4];
wire w_pp_31_05 = i_multiplier[31] & i_multiplicand[ 5];
wire w_pp_31_06 = i_multiplier[31] & i_multiplicand[ 6];
wire w_pp_31_07 = i_multiplier[31] & i_multiplicand[ 7];
wire w_pp_31_08 = i_multiplier[31] & i_multiplicand[ 8];
wire w_pp_31_09 = i_multiplier[31] & i_multiplicand[ 9];
wire w_pp_31_10 = i_multiplier[31] & i_multiplicand[10];
wire w_pp_31_11 = i_multiplier[31] & i_multiplicand[11];
wire w_pp_31_12 = i_multiplier[31] & i_multiplicand[12];
wire w_pp_31_13 = i_multiplier[31] & i_multiplicand[13];
wire w_pp_31_14 = i_multiplier[31] & i_multiplicand[14];
wire w_pp_31_15 = i_multiplier[31] & i_multiplicand[15];
wire w_pp_31_16 = i_multiplier[31] & i_multiplicand[16];
wire w_pp_31_17 = i_multiplier[31] & i_multiplicand[17];
wire w_pp_31_18 = i_multiplier[31] & i_multiplicand[18];
wire w_pp_31_19 = i_multiplier[31] & i_multiplicand[19];
wire w_pp_31_20 = i_multiplier[31] & i_multiplicand[20];
wire w_pp_31_21 = i_multiplier[31] & i_multiplicand[21];
wire w_pp_31_22 = i_multiplier[31] & i_multiplicand[22];
wire w_pp_31_23 = i_multiplier[31] & i_multiplicand[23];
wire w_pp_31_24 = i_multiplier[31] & i_multiplicand[24];
wire w_pp_31_25 = i_multiplier[31] & i_multiplicand[25];
wire w_pp_31_26 = i_multiplier[31] & i_multiplicand[26];
wire w_pp_31_27 = i_multiplier[31] & i_multiplicand[27];
wire w_pp_31_28 = i_multiplier[31] & i_multiplicand[28];
wire w_pp_31_29 = i_multiplier[31] & i_multiplicand[29];
wire w_pp_31_30 = i_multiplier[31] & i_multiplicand[30];
wire w_pp_31_31 = i_multiplier[31] & i_multiplicand[31];

// Partial products reduction using Wallace tree
wire w_sum_01_02, w_carry_01_02;
math_adder_half HA_01_02(.i_a(w_pp_00_01), .i_b(w_pp_01_00), .ow_sum(w_sum_01_02), .ow_carry(w_carry_01_02));
wire w_sum_02_04, w_carry_02_04;
math_adder_full FA_02_04(.i_a(w_pp_00_02), .i_b(w_pp_01_01), .i_c(w_pp_02_00), .ow_sum(w_sum_02_04), .ow_carry(w_carry_02_04));
wire w_sum_02_02, w_carry_02_02;
math_adder_half HA_02_02(.i_a(w_carry_01_02), .i_b(w_sum_02_04), .ow_sum(w_sum_02_02), .ow_carry(w_carry_02_02));
wire w_sum_03_06, w_carry_03_06;
math_adder_full FA_03_06(.i_a(w_pp_00_03), .i_b(w_pp_01_02), .i_c(w_pp_02_01), .ow_sum(w_sum_03_06), .ow_carry(w_carry_03_06));
wire w_sum_03_04, w_carry_03_04;
math_adder_full FA_03_04(.i_a(w_pp_03_00), .i_b(w_carry_02_04), .i_c(w_carry_02_02), .ow_sum(w_sum_03_04), .ow_carry(w_carry_03_04));
wire w_sum_03_02, w_carry_03_02;
math_adder_half HA_03_02(.i_a(w_sum_03_06), .i_b(w_sum_03_04), .ow_sum(w_sum_03_02), .ow_carry(w_carry_03_02));
wire w_sum_04_08, w_carry_04_08;
math_adder_full FA_04_08(.i_a(w_pp_00_04), .i_b(w_pp_01_03), .i_c(w_pp_02_02), .ow_sum(w_sum_04_08), .ow_carry(w_carry_04_08));
wire w_sum_04_06, w_carry_04_06;
math_adder_full FA_04_06(.i_a(w_pp_03_01), .i_b(w_pp_04_00), .i_c(w_carry_03_06), .ow_sum(w_sum_04_06), .ow_carry(w_carry_04_06));
wire w_sum_04_04, w_carry_04_04;
math_adder_full FA_04_04(.i_a(w_carry_03_04), .i_b(w_carry_03_02), .i_c(w_sum_04_08), .ow_sum(w_sum_04_04), .ow_carry(w_carry_04_04));
wire w_sum_04_02, w_carry_04_02;
math_adder_half HA_04_02(.i_a(w_sum_04_06), .i_b(w_sum_04_04), .ow_sum(w_sum_04_02), .ow_carry(w_carry_04_02));
wire w_sum_05_10, w_carry_05_10;
math_adder_full FA_05_10(.i_a(w_pp_00_05), .i_b(w_pp_01_04), .i_c(w_pp_02_03), .ow_sum(w_sum_05_10), .ow_carry(w_carry_05_10));
wire w_sum_05_08, w_carry_05_08;
math_adder_full FA_05_08(.i_a(w_pp_03_02), .i_b(w_pp_04_01), .i_c(w_pp_05_00), .ow_sum(w_sum_05_08), .ow_carry(w_carry_05_08));
wire w_sum_05_06, w_carry_05_06;
math_adder_full FA_05_06(.i_a(w_carry_04_08), .i_b(w_carry_04_06), .i_c(w_carry_04_04), .ow_sum(w_sum_05_06), .ow_carry(w_carry_05_06));
wire w_sum_05_04, w_carry_05_04;
math_adder_full FA_05_04(.i_a(w_carry_04_02), .i_b(w_sum_05_10), .i_c(w_sum_05_08), .ow_sum(w_sum_05_04), .ow_carry(w_carry_05_04));
wire w_sum_05_02, w_carry_05_02;
math_adder_half HA_05_02(.i_a(w_sum_05_06), .i_b(w_sum_05_04), .ow_sum(w_sum_05_02), .ow_carry(w_carry_05_02));
wire w_sum_06_12, w_carry_06_12;
math_adder_full FA_06_12(.i_a(w_pp_00_06), .i_b(w_pp_01_05), .i_c(w_pp_02_04), .ow_sum(w_sum_06_12), .ow_carry(w_carry_06_12));
wire w_sum_06_10, w_carry_06_10;
math_adder_full FA_06_10(.i_a(w_pp_03_03), .i_b(w_pp_04_02), .i_c(w_pp_05_01), .ow_sum(w_sum_06_10), .ow_carry(w_carry_06_10));
wire w_sum_06_08, w_carry_06_08;
math_adder_full FA_06_08(.i_a(w_pp_06_00), .i_b(w_carry_05_10), .i_c(w_carry_05_08), .ow_sum(w_sum_06_08), .ow_carry(w_carry_06_08));
wire w_sum_06_06, w_carry_06_06;
math_adder_full FA_06_06(.i_a(w_carry_05_06), .i_b(w_carry_05_04), .i_c(w_carry_05_02), .ow_sum(w_sum_06_06), .ow_carry(w_carry_06_06));
wire w_sum_06_04, w_carry_06_04;
math_adder_full FA_06_04(.i_a(w_sum_06_12), .i_b(w_sum_06_10), .i_c(w_sum_06_08), .ow_sum(w_sum_06_04), .ow_carry(w_carry_06_04));
wire w_sum_06_02, w_carry_06_02;
math_adder_half HA_06_02(.i_a(w_sum_06_06), .i_b(w_sum_06_04), .ow_sum(w_sum_06_02), .ow_carry(w_carry_06_02));
wire w_sum_07_14, w_carry_07_14;
math_adder_full FA_07_14(.i_a(w_pp_00_07), .i_b(w_pp_01_06), .i_c(w_pp_02_05), .ow_sum(w_sum_07_14), .ow_carry(w_carry_07_14));
wire w_sum_07_12, w_carry_07_12;
math_adder_full FA_07_12(.i_a(w_pp_03_04), .i_b(w_pp_04_03), .i_c(w_pp_05_02), .ow_sum(w_sum_07_12), .ow_carry(w_carry_07_12));
wire w_sum_07_10, w_carry_07_10;
math_adder_full FA_07_10(.i_a(w_pp_06_01), .i_b(w_pp_07_00), .i_c(w_carry_06_12), .ow_sum(w_sum_07_10), .ow_carry(w_carry_07_10));
wire w_sum_07_08, w_carry_07_08;
math_adder_full FA_07_08(.i_a(w_carry_06_10), .i_b(w_carry_06_08), .i_c(w_carry_06_06), .ow_sum(w_sum_07_08), .ow_carry(w_carry_07_08));
wire w_sum_07_06, w_carry_07_06;
math_adder_full FA_07_06(.i_a(w_carry_06_04), .i_b(w_carry_06_02), .i_c(w_sum_07_14), .ow_sum(w_sum_07_06), .ow_carry(w_carry_07_06));
wire w_sum_07_04, w_carry_07_04;
math_adder_full FA_07_04(.i_a(w_sum_07_12), .i_b(w_sum_07_10), .i_c(w_sum_07_08), .ow_sum(w_sum_07_04), .ow_carry(w_carry_07_04));
wire w_sum_07_02, w_carry_07_02;
math_adder_half HA_07_02(.i_a(w_sum_07_06), .i_b(w_sum_07_04), .ow_sum(w_sum_07_02), .ow_carry(w_carry_07_02));
wire w_sum_08_16, w_carry_08_16;
math_adder_full FA_08_16(.i_a(w_pp_00_08), .i_b(w_pp_01_07), .i_c(w_pp_02_06), .ow_sum(w_sum_08_16), .ow_carry(w_carry_08_16));
wire w_sum_08_14, w_carry_08_14;
math_adder_full FA_08_14(.i_a(w_pp_03_05), .i_b(w_pp_04_04), .i_c(w_pp_05_03), .ow_sum(w_sum_08_14), .ow_carry(w_carry_08_14));
wire w_sum_08_12, w_carry_08_12;
math_adder_full FA_08_12(.i_a(w_pp_06_02), .i_b(w_pp_07_01), .i_c(w_pp_08_00), .ow_sum(w_sum_08_12), .ow_carry(w_carry_08_12));
wire w_sum_08_10, w_carry_08_10;
math_adder_full FA_08_10(.i_a(w_carry_07_14), .i_b(w_carry_07_12), .i_c(w_carry_07_10), .ow_sum(w_sum_08_10), .ow_carry(w_carry_08_10));
wire w_sum_08_08, w_carry_08_08;
math_adder_full FA_08_08(.i_a(w_carry_07_08), .i_b(w_carry_07_06), .i_c(w_carry_07_04), .ow_sum(w_sum_08_08), .ow_carry(w_carry_08_08));
wire w_sum_08_06, w_carry_08_06;
math_adder_full FA_08_06(.i_a(w_carry_07_02), .i_b(w_sum_08_16), .i_c(w_sum_08_14), .ow_sum(w_sum_08_06), .ow_carry(w_carry_08_06));
wire w_sum_08_04, w_carry_08_04;
math_adder_full FA_08_04(.i_a(w_sum_08_12), .i_b(w_sum_08_10), .i_c(w_sum_08_08), .ow_sum(w_sum_08_04), .ow_carry(w_carry_08_04));
wire w_sum_08_02, w_carry_08_02;
math_adder_half HA_08_02(.i_a(w_sum_08_06), .i_b(w_sum_08_04), .ow_sum(w_sum_08_02), .ow_carry(w_carry_08_02));
wire w_sum_09_18, w_carry_09_18;
math_adder_full FA_09_18(.i_a(w_pp_00_09), .i_b(w_pp_01_08), .i_c(w_pp_02_07), .ow_sum(w_sum_09_18), .ow_carry(w_carry_09_18));
wire w_sum_09_16, w_carry_09_16;
math_adder_full FA_09_16(.i_a(w_pp_03_06), .i_b(w_pp_04_05), .i_c(w_pp_05_04), .ow_sum(w_sum_09_16), .ow_carry(w_carry_09_16));
wire w_sum_09_14, w_carry_09_14;
math_adder_full FA_09_14(.i_a(w_pp_06_03), .i_b(w_pp_07_02), .i_c(w_pp_08_01), .ow_sum(w_sum_09_14), .ow_carry(w_carry_09_14));
wire w_sum_09_12, w_carry_09_12;
math_adder_full FA_09_12(.i_a(w_pp_09_00), .i_b(w_carry_08_16), .i_c(w_carry_08_14), .ow_sum(w_sum_09_12), .ow_carry(w_carry_09_12));
wire w_sum_09_10, w_carry_09_10;
math_adder_full FA_09_10(.i_a(w_carry_08_12), .i_b(w_carry_08_10), .i_c(w_carry_08_08), .ow_sum(w_sum_09_10), .ow_carry(w_carry_09_10));
wire w_sum_09_08, w_carry_09_08;
math_adder_full FA_09_08(.i_a(w_carry_08_06), .i_b(w_carry_08_04), .i_c(w_carry_08_02), .ow_sum(w_sum_09_08), .ow_carry(w_carry_09_08));
wire w_sum_09_06, w_carry_09_06;
math_adder_full FA_09_06(.i_a(w_sum_09_18), .i_b(w_sum_09_16), .i_c(w_sum_09_14), .ow_sum(w_sum_09_06), .ow_carry(w_carry_09_06));
wire w_sum_09_04, w_carry_09_04;
math_adder_full FA_09_04(.i_a(w_sum_09_12), .i_b(w_sum_09_10), .i_c(w_sum_09_08), .ow_sum(w_sum_09_04), .ow_carry(w_carry_09_04));
wire w_sum_09_02, w_carry_09_02;
math_adder_half HA_09_02(.i_a(w_sum_09_06), .i_b(w_sum_09_04), .ow_sum(w_sum_09_02), .ow_carry(w_carry_09_02));
wire w_sum_10_20, w_carry_10_20;
math_adder_full FA_10_20(.i_a(w_pp_00_10), .i_b(w_pp_01_09), .i_c(w_pp_02_08), .ow_sum(w_sum_10_20), .ow_carry(w_carry_10_20));
wire w_sum_10_18, w_carry_10_18;
math_adder_full FA_10_18(.i_a(w_pp_03_07), .i_b(w_pp_04_06), .i_c(w_pp_05_05), .ow_sum(w_sum_10_18), .ow_carry(w_carry_10_18));
wire w_sum_10_16, w_carry_10_16;
math_adder_full FA_10_16(.i_a(w_pp_06_04), .i_b(w_pp_07_03), .i_c(w_pp_08_02), .ow_sum(w_sum_10_16), .ow_carry(w_carry_10_16));
wire w_sum_10_14, w_carry_10_14;
math_adder_full FA_10_14(.i_a(w_pp_09_01), .i_b(w_pp_10_00), .i_c(w_carry_09_18), .ow_sum(w_sum_10_14), .ow_carry(w_carry_10_14));
wire w_sum_10_12, w_carry_10_12;
math_adder_full FA_10_12(.i_a(w_carry_09_16), .i_b(w_carry_09_14), .i_c(w_carry_09_12), .ow_sum(w_sum_10_12), .ow_carry(w_carry_10_12));
wire w_sum_10_10, w_carry_10_10;
math_adder_full FA_10_10(.i_a(w_carry_09_10), .i_b(w_carry_09_08), .i_c(w_carry_09_06), .ow_sum(w_sum_10_10), .ow_carry(w_carry_10_10));
wire w_sum_10_08, w_carry_10_08;
math_adder_full FA_10_08(.i_a(w_carry_09_04), .i_b(w_carry_09_02), .i_c(w_sum_10_20), .ow_sum(w_sum_10_08), .ow_carry(w_carry_10_08));
wire w_sum_10_06, w_carry_10_06;
math_adder_full FA_10_06(.i_a(w_sum_10_18), .i_b(w_sum_10_16), .i_c(w_sum_10_14), .ow_sum(w_sum_10_06), .ow_carry(w_carry_10_06));
wire w_sum_10_04, w_carry_10_04;
math_adder_full FA_10_04(.i_a(w_sum_10_12), .i_b(w_sum_10_10), .i_c(w_sum_10_08), .ow_sum(w_sum_10_04), .ow_carry(w_carry_10_04));
wire w_sum_10_02, w_carry_10_02;
math_adder_half HA_10_02(.i_a(w_sum_10_06), .i_b(w_sum_10_04), .ow_sum(w_sum_10_02), .ow_carry(w_carry_10_02));
wire w_sum_11_22, w_carry_11_22;
math_adder_full FA_11_22(.i_a(w_pp_00_11), .i_b(w_pp_01_10), .i_c(w_pp_02_09), .ow_sum(w_sum_11_22), .ow_carry(w_carry_11_22));
wire w_sum_11_20, w_carry_11_20;
math_adder_full FA_11_20(.i_a(w_pp_03_08), .i_b(w_pp_04_07), .i_c(w_pp_05_06), .ow_sum(w_sum_11_20), .ow_carry(w_carry_11_20));
wire w_sum_11_18, w_carry_11_18;
math_adder_full FA_11_18(.i_a(w_pp_06_05), .i_b(w_pp_07_04), .i_c(w_pp_08_03), .ow_sum(w_sum_11_18), .ow_carry(w_carry_11_18));
wire w_sum_11_16, w_carry_11_16;
math_adder_full FA_11_16(.i_a(w_pp_09_02), .i_b(w_pp_10_01), .i_c(w_pp_11_00), .ow_sum(w_sum_11_16), .ow_carry(w_carry_11_16));
wire w_sum_11_14, w_carry_11_14;
math_adder_full FA_11_14(.i_a(w_carry_10_20), .i_b(w_carry_10_18), .i_c(w_carry_10_16), .ow_sum(w_sum_11_14), .ow_carry(w_carry_11_14));
wire w_sum_11_12, w_carry_11_12;
math_adder_full FA_11_12(.i_a(w_carry_10_14), .i_b(w_carry_10_12), .i_c(w_carry_10_10), .ow_sum(w_sum_11_12), .ow_carry(w_carry_11_12));
wire w_sum_11_10, w_carry_11_10;
math_adder_full FA_11_10(.i_a(w_carry_10_08), .i_b(w_carry_10_06), .i_c(w_carry_10_04), .ow_sum(w_sum_11_10), .ow_carry(w_carry_11_10));
wire w_sum_11_08, w_carry_11_08;
math_adder_full FA_11_08(.i_a(w_carry_10_02), .i_b(w_sum_11_22), .i_c(w_sum_11_20), .ow_sum(w_sum_11_08), .ow_carry(w_carry_11_08));
wire w_sum_11_06, w_carry_11_06;
math_adder_full FA_11_06(.i_a(w_sum_11_18), .i_b(w_sum_11_16), .i_c(w_sum_11_14), .ow_sum(w_sum_11_06), .ow_carry(w_carry_11_06));
wire w_sum_11_04, w_carry_11_04;
math_adder_full FA_11_04(.i_a(w_sum_11_12), .i_b(w_sum_11_10), .i_c(w_sum_11_08), .ow_sum(w_sum_11_04), .ow_carry(w_carry_11_04));
wire w_sum_11_02, w_carry_11_02;
math_adder_half HA_11_02(.i_a(w_sum_11_06), .i_b(w_sum_11_04), .ow_sum(w_sum_11_02), .ow_carry(w_carry_11_02));
wire w_sum_12_24, w_carry_12_24;
math_adder_full FA_12_24(.i_a(w_pp_00_12), .i_b(w_pp_01_11), .i_c(w_pp_02_10), .ow_sum(w_sum_12_24), .ow_carry(w_carry_12_24));
wire w_sum_12_22, w_carry_12_22;
math_adder_full FA_12_22(.i_a(w_pp_03_09), .i_b(w_pp_04_08), .i_c(w_pp_05_07), .ow_sum(w_sum_12_22), .ow_carry(w_carry_12_22));
wire w_sum_12_20, w_carry_12_20;
math_adder_full FA_12_20(.i_a(w_pp_06_06), .i_b(w_pp_07_05), .i_c(w_pp_08_04), .ow_sum(w_sum_12_20), .ow_carry(w_carry_12_20));
wire w_sum_12_18, w_carry_12_18;
math_adder_full FA_12_18(.i_a(w_pp_09_03), .i_b(w_pp_10_02), .i_c(w_pp_11_01), .ow_sum(w_sum_12_18), .ow_carry(w_carry_12_18));
wire w_sum_12_16, w_carry_12_16;
math_adder_full FA_12_16(.i_a(w_pp_12_00), .i_b(w_carry_11_22), .i_c(w_carry_11_20), .ow_sum(w_sum_12_16), .ow_carry(w_carry_12_16));
wire w_sum_12_14, w_carry_12_14;
math_adder_full FA_12_14(.i_a(w_carry_11_18), .i_b(w_carry_11_16), .i_c(w_carry_11_14), .ow_sum(w_sum_12_14), .ow_carry(w_carry_12_14));
wire w_sum_12_12, w_carry_12_12;
math_adder_full FA_12_12(.i_a(w_carry_11_12), .i_b(w_carry_11_10), .i_c(w_carry_11_08), .ow_sum(w_sum_12_12), .ow_carry(w_carry_12_12));
wire w_sum_12_10, w_carry_12_10;
math_adder_full FA_12_10(.i_a(w_carry_11_06), .i_b(w_carry_11_04), .i_c(w_carry_11_02), .ow_sum(w_sum_12_10), .ow_carry(w_carry_12_10));
wire w_sum_12_08, w_carry_12_08;
math_adder_full FA_12_08(.i_a(w_sum_12_24), .i_b(w_sum_12_22), .i_c(w_sum_12_20), .ow_sum(w_sum_12_08), .ow_carry(w_carry_12_08));
wire w_sum_12_06, w_carry_12_06;
math_adder_full FA_12_06(.i_a(w_sum_12_18), .i_b(w_sum_12_16), .i_c(w_sum_12_14), .ow_sum(w_sum_12_06), .ow_carry(w_carry_12_06));
wire w_sum_12_04, w_carry_12_04;
math_adder_full FA_12_04(.i_a(w_sum_12_12), .i_b(w_sum_12_10), .i_c(w_sum_12_08), .ow_sum(w_sum_12_04), .ow_carry(w_carry_12_04));
wire w_sum_12_02, w_carry_12_02;
math_adder_half HA_12_02(.i_a(w_sum_12_06), .i_b(w_sum_12_04), .ow_sum(w_sum_12_02), .ow_carry(w_carry_12_02));
wire w_sum_13_26, w_carry_13_26;
math_adder_full FA_13_26(.i_a(w_pp_00_13), .i_b(w_pp_01_12), .i_c(w_pp_02_11), .ow_sum(w_sum_13_26), .ow_carry(w_carry_13_26));
wire w_sum_13_24, w_carry_13_24;
math_adder_full FA_13_24(.i_a(w_pp_03_10), .i_b(w_pp_04_09), .i_c(w_pp_05_08), .ow_sum(w_sum_13_24), .ow_carry(w_carry_13_24));
wire w_sum_13_22, w_carry_13_22;
math_adder_full FA_13_22(.i_a(w_pp_06_07), .i_b(w_pp_07_06), .i_c(w_pp_08_05), .ow_sum(w_sum_13_22), .ow_carry(w_carry_13_22));
wire w_sum_13_20, w_carry_13_20;
math_adder_full FA_13_20(.i_a(w_pp_09_04), .i_b(w_pp_10_03), .i_c(w_pp_11_02), .ow_sum(w_sum_13_20), .ow_carry(w_carry_13_20));
wire w_sum_13_18, w_carry_13_18;
math_adder_full FA_13_18(.i_a(w_pp_12_01), .i_b(w_pp_13_00), .i_c(w_carry_12_24), .ow_sum(w_sum_13_18), .ow_carry(w_carry_13_18));
wire w_sum_13_16, w_carry_13_16;
math_adder_full FA_13_16(.i_a(w_carry_12_22), .i_b(w_carry_12_20), .i_c(w_carry_12_18), .ow_sum(w_sum_13_16), .ow_carry(w_carry_13_16));
wire w_sum_13_14, w_carry_13_14;
math_adder_full FA_13_14(.i_a(w_carry_12_16), .i_b(w_carry_12_14), .i_c(w_carry_12_12), .ow_sum(w_sum_13_14), .ow_carry(w_carry_13_14));
wire w_sum_13_12, w_carry_13_12;
math_adder_full FA_13_12(.i_a(w_carry_12_10), .i_b(w_carry_12_08), .i_c(w_carry_12_06), .ow_sum(w_sum_13_12), .ow_carry(w_carry_13_12));
wire w_sum_13_10, w_carry_13_10;
math_adder_full FA_13_10(.i_a(w_carry_12_04), .i_b(w_carry_12_02), .i_c(w_sum_13_26), .ow_sum(w_sum_13_10), .ow_carry(w_carry_13_10));
wire w_sum_13_08, w_carry_13_08;
math_adder_full FA_13_08(.i_a(w_sum_13_24), .i_b(w_sum_13_22), .i_c(w_sum_13_20), .ow_sum(w_sum_13_08), .ow_carry(w_carry_13_08));
wire w_sum_13_06, w_carry_13_06;
math_adder_full FA_13_06(.i_a(w_sum_13_18), .i_b(w_sum_13_16), .i_c(w_sum_13_14), .ow_sum(w_sum_13_06), .ow_carry(w_carry_13_06));
wire w_sum_13_04, w_carry_13_04;
math_adder_full FA_13_04(.i_a(w_sum_13_12), .i_b(w_sum_13_10), .i_c(w_sum_13_08), .ow_sum(w_sum_13_04), .ow_carry(w_carry_13_04));
wire w_sum_13_02, w_carry_13_02;
math_adder_half HA_13_02(.i_a(w_sum_13_06), .i_b(w_sum_13_04), .ow_sum(w_sum_13_02), .ow_carry(w_carry_13_02));
wire w_sum_14_28, w_carry_14_28;
math_adder_full FA_14_28(.i_a(w_pp_00_14), .i_b(w_pp_01_13), .i_c(w_pp_02_12), .ow_sum(w_sum_14_28), .ow_carry(w_carry_14_28));
wire w_sum_14_26, w_carry_14_26;
math_adder_full FA_14_26(.i_a(w_pp_03_11), .i_b(w_pp_04_10), .i_c(w_pp_05_09), .ow_sum(w_sum_14_26), .ow_carry(w_carry_14_26));
wire w_sum_14_24, w_carry_14_24;
math_adder_full FA_14_24(.i_a(w_pp_06_08), .i_b(w_pp_07_07), .i_c(w_pp_08_06), .ow_sum(w_sum_14_24), .ow_carry(w_carry_14_24));
wire w_sum_14_22, w_carry_14_22;
math_adder_full FA_14_22(.i_a(w_pp_09_05), .i_b(w_pp_10_04), .i_c(w_pp_11_03), .ow_sum(w_sum_14_22), .ow_carry(w_carry_14_22));
wire w_sum_14_20, w_carry_14_20;
math_adder_full FA_14_20(.i_a(w_pp_12_02), .i_b(w_pp_13_01), .i_c(w_pp_14_00), .ow_sum(w_sum_14_20), .ow_carry(w_carry_14_20));
wire w_sum_14_18, w_carry_14_18;
math_adder_full FA_14_18(.i_a(w_carry_13_26), .i_b(w_carry_13_24), .i_c(w_carry_13_22), .ow_sum(w_sum_14_18), .ow_carry(w_carry_14_18));
wire w_sum_14_16, w_carry_14_16;
math_adder_full FA_14_16(.i_a(w_carry_13_20), .i_b(w_carry_13_18), .i_c(w_carry_13_16), .ow_sum(w_sum_14_16), .ow_carry(w_carry_14_16));
wire w_sum_14_14, w_carry_14_14;
math_adder_full FA_14_14(.i_a(w_carry_13_14), .i_b(w_carry_13_12), .i_c(w_carry_13_10), .ow_sum(w_sum_14_14), .ow_carry(w_carry_14_14));
wire w_sum_14_12, w_carry_14_12;
math_adder_full FA_14_12(.i_a(w_carry_13_08), .i_b(w_carry_13_06), .i_c(w_carry_13_04), .ow_sum(w_sum_14_12), .ow_carry(w_carry_14_12));
wire w_sum_14_10, w_carry_14_10;
math_adder_full FA_14_10(.i_a(w_carry_13_02), .i_b(w_sum_14_28), .i_c(w_sum_14_26), .ow_sum(w_sum_14_10), .ow_carry(w_carry_14_10));
wire w_sum_14_08, w_carry_14_08;
math_adder_full FA_14_08(.i_a(w_sum_14_24), .i_b(w_sum_14_22), .i_c(w_sum_14_20), .ow_sum(w_sum_14_08), .ow_carry(w_carry_14_08));
wire w_sum_14_06, w_carry_14_06;
math_adder_full FA_14_06(.i_a(w_sum_14_18), .i_b(w_sum_14_16), .i_c(w_sum_14_14), .ow_sum(w_sum_14_06), .ow_carry(w_carry_14_06));
wire w_sum_14_04, w_carry_14_04;
math_adder_full FA_14_04(.i_a(w_sum_14_12), .i_b(w_sum_14_10), .i_c(w_sum_14_08), .ow_sum(w_sum_14_04), .ow_carry(w_carry_14_04));
wire w_sum_14_02, w_carry_14_02;
math_adder_half HA_14_02(.i_a(w_sum_14_06), .i_b(w_sum_14_04), .ow_sum(w_sum_14_02), .ow_carry(w_carry_14_02));
wire w_sum_15_30, w_carry_15_30;
math_adder_full FA_15_30(.i_a(w_pp_00_15), .i_b(w_pp_01_14), .i_c(w_pp_02_13), .ow_sum(w_sum_15_30), .ow_carry(w_carry_15_30));
wire w_sum_15_28, w_carry_15_28;
math_adder_full FA_15_28(.i_a(w_pp_03_12), .i_b(w_pp_04_11), .i_c(w_pp_05_10), .ow_sum(w_sum_15_28), .ow_carry(w_carry_15_28));
wire w_sum_15_26, w_carry_15_26;
math_adder_full FA_15_26(.i_a(w_pp_06_09), .i_b(w_pp_07_08), .i_c(w_pp_08_07), .ow_sum(w_sum_15_26), .ow_carry(w_carry_15_26));
wire w_sum_15_24, w_carry_15_24;
math_adder_full FA_15_24(.i_a(w_pp_09_06), .i_b(w_pp_10_05), .i_c(w_pp_11_04), .ow_sum(w_sum_15_24), .ow_carry(w_carry_15_24));
wire w_sum_15_22, w_carry_15_22;
math_adder_full FA_15_22(.i_a(w_pp_12_03), .i_b(w_pp_13_02), .i_c(w_pp_14_01), .ow_sum(w_sum_15_22), .ow_carry(w_carry_15_22));
wire w_sum_15_20, w_carry_15_20;
math_adder_full FA_15_20(.i_a(w_pp_15_00), .i_b(w_carry_14_28), .i_c(w_carry_14_26), .ow_sum(w_sum_15_20), .ow_carry(w_carry_15_20));
wire w_sum_15_18, w_carry_15_18;
math_adder_full FA_15_18(.i_a(w_carry_14_24), .i_b(w_carry_14_22), .i_c(w_carry_14_20), .ow_sum(w_sum_15_18), .ow_carry(w_carry_15_18));
wire w_sum_15_16, w_carry_15_16;
math_adder_full FA_15_16(.i_a(w_carry_14_18), .i_b(w_carry_14_16), .i_c(w_carry_14_14), .ow_sum(w_sum_15_16), .ow_carry(w_carry_15_16));
wire w_sum_15_14, w_carry_15_14;
math_adder_full FA_15_14(.i_a(w_carry_14_12), .i_b(w_carry_14_10), .i_c(w_carry_14_08), .ow_sum(w_sum_15_14), .ow_carry(w_carry_15_14));
wire w_sum_15_12, w_carry_15_12;
math_adder_full FA_15_12(.i_a(w_carry_14_06), .i_b(w_carry_14_04), .i_c(w_carry_14_02), .ow_sum(w_sum_15_12), .ow_carry(w_carry_15_12));
wire w_sum_15_10, w_carry_15_10;
math_adder_full FA_15_10(.i_a(w_sum_15_30), .i_b(w_sum_15_28), .i_c(w_sum_15_26), .ow_sum(w_sum_15_10), .ow_carry(w_carry_15_10));
wire w_sum_15_08, w_carry_15_08;
math_adder_full FA_15_08(.i_a(w_sum_15_24), .i_b(w_sum_15_22), .i_c(w_sum_15_20), .ow_sum(w_sum_15_08), .ow_carry(w_carry_15_08));
wire w_sum_15_06, w_carry_15_06;
math_adder_full FA_15_06(.i_a(w_sum_15_18), .i_b(w_sum_15_16), .i_c(w_sum_15_14), .ow_sum(w_sum_15_06), .ow_carry(w_carry_15_06));
wire w_sum_15_04, w_carry_15_04;
math_adder_full FA_15_04(.i_a(w_sum_15_12), .i_b(w_sum_15_10), .i_c(w_sum_15_08), .ow_sum(w_sum_15_04), .ow_carry(w_carry_15_04));
wire w_sum_15_02, w_carry_15_02;
math_adder_half HA_15_02(.i_a(w_sum_15_06), .i_b(w_sum_15_04), .ow_sum(w_sum_15_02), .ow_carry(w_carry_15_02));
wire w_sum_16_32, w_carry_16_32;
math_adder_full FA_16_32(.i_a(w_pp_00_16), .i_b(w_pp_01_15), .i_c(w_pp_02_14), .ow_sum(w_sum_16_32), .ow_carry(w_carry_16_32));
wire w_sum_16_30, w_carry_16_30;
math_adder_full FA_16_30(.i_a(w_pp_03_13), .i_b(w_pp_04_12), .i_c(w_pp_05_11), .ow_sum(w_sum_16_30), .ow_carry(w_carry_16_30));
wire w_sum_16_28, w_carry_16_28;
math_adder_full FA_16_28(.i_a(w_pp_06_10), .i_b(w_pp_07_09), .i_c(w_pp_08_08), .ow_sum(w_sum_16_28), .ow_carry(w_carry_16_28));
wire w_sum_16_26, w_carry_16_26;
math_adder_full FA_16_26(.i_a(w_pp_09_07), .i_b(w_pp_10_06), .i_c(w_pp_11_05), .ow_sum(w_sum_16_26), .ow_carry(w_carry_16_26));
wire w_sum_16_24, w_carry_16_24;
math_adder_full FA_16_24(.i_a(w_pp_12_04), .i_b(w_pp_13_03), .i_c(w_pp_14_02), .ow_sum(w_sum_16_24), .ow_carry(w_carry_16_24));
wire w_sum_16_22, w_carry_16_22;
math_adder_full FA_16_22(.i_a(w_pp_15_01), .i_b(w_pp_16_00), .i_c(w_carry_15_30), .ow_sum(w_sum_16_22), .ow_carry(w_carry_16_22));
wire w_sum_16_20, w_carry_16_20;
math_adder_full FA_16_20(.i_a(w_carry_15_28), .i_b(w_carry_15_26), .i_c(w_carry_15_24), .ow_sum(w_sum_16_20), .ow_carry(w_carry_16_20));
wire w_sum_16_18, w_carry_16_18;
math_adder_full FA_16_18(.i_a(w_carry_15_22), .i_b(w_carry_15_20), .i_c(w_carry_15_18), .ow_sum(w_sum_16_18), .ow_carry(w_carry_16_18));
wire w_sum_16_16, w_carry_16_16;
math_adder_full FA_16_16(.i_a(w_carry_15_16), .i_b(w_carry_15_14), .i_c(w_carry_15_12), .ow_sum(w_sum_16_16), .ow_carry(w_carry_16_16));
wire w_sum_16_14, w_carry_16_14;
math_adder_full FA_16_14(.i_a(w_carry_15_10), .i_b(w_carry_15_08), .i_c(w_carry_15_06), .ow_sum(w_sum_16_14), .ow_carry(w_carry_16_14));
wire w_sum_16_12, w_carry_16_12;
math_adder_full FA_16_12(.i_a(w_carry_15_04), .i_b(w_carry_15_02), .i_c(w_sum_16_32), .ow_sum(w_sum_16_12), .ow_carry(w_carry_16_12));
wire w_sum_16_10, w_carry_16_10;
math_adder_full FA_16_10(.i_a(w_sum_16_30), .i_b(w_sum_16_28), .i_c(w_sum_16_26), .ow_sum(w_sum_16_10), .ow_carry(w_carry_16_10));
wire w_sum_16_08, w_carry_16_08;
math_adder_full FA_16_08(.i_a(w_sum_16_24), .i_b(w_sum_16_22), .i_c(w_sum_16_20), .ow_sum(w_sum_16_08), .ow_carry(w_carry_16_08));
wire w_sum_16_06, w_carry_16_06;
math_adder_full FA_16_06(.i_a(w_sum_16_18), .i_b(w_sum_16_16), .i_c(w_sum_16_14), .ow_sum(w_sum_16_06), .ow_carry(w_carry_16_06));
wire w_sum_16_04, w_carry_16_04;
math_adder_full FA_16_04(.i_a(w_sum_16_12), .i_b(w_sum_16_10), .i_c(w_sum_16_08), .ow_sum(w_sum_16_04), .ow_carry(w_carry_16_04));
wire w_sum_16_02, w_carry_16_02;
math_adder_half HA_16_02(.i_a(w_sum_16_06), .i_b(w_sum_16_04), .ow_sum(w_sum_16_02), .ow_carry(w_carry_16_02));
wire w_sum_17_34, w_carry_17_34;
math_adder_full FA_17_34(.i_a(w_pp_00_17), .i_b(w_pp_01_16), .i_c(w_pp_02_15), .ow_sum(w_sum_17_34), .ow_carry(w_carry_17_34));
wire w_sum_17_32, w_carry_17_32;
math_adder_full FA_17_32(.i_a(w_pp_03_14), .i_b(w_pp_04_13), .i_c(w_pp_05_12), .ow_sum(w_sum_17_32), .ow_carry(w_carry_17_32));
wire w_sum_17_30, w_carry_17_30;
math_adder_full FA_17_30(.i_a(w_pp_06_11), .i_b(w_pp_07_10), .i_c(w_pp_08_09), .ow_sum(w_sum_17_30), .ow_carry(w_carry_17_30));
wire w_sum_17_28, w_carry_17_28;
math_adder_full FA_17_28(.i_a(w_pp_09_08), .i_b(w_pp_10_07), .i_c(w_pp_11_06), .ow_sum(w_sum_17_28), .ow_carry(w_carry_17_28));
wire w_sum_17_26, w_carry_17_26;
math_adder_full FA_17_26(.i_a(w_pp_12_05), .i_b(w_pp_13_04), .i_c(w_pp_14_03), .ow_sum(w_sum_17_26), .ow_carry(w_carry_17_26));
wire w_sum_17_24, w_carry_17_24;
math_adder_full FA_17_24(.i_a(w_pp_15_02), .i_b(w_pp_16_01), .i_c(w_pp_17_00), .ow_sum(w_sum_17_24), .ow_carry(w_carry_17_24));
wire w_sum_17_22, w_carry_17_22;
math_adder_full FA_17_22(.i_a(w_carry_16_32), .i_b(w_carry_16_30), .i_c(w_carry_16_28), .ow_sum(w_sum_17_22), .ow_carry(w_carry_17_22));
wire w_sum_17_20, w_carry_17_20;
math_adder_full FA_17_20(.i_a(w_carry_16_26), .i_b(w_carry_16_24), .i_c(w_carry_16_22), .ow_sum(w_sum_17_20), .ow_carry(w_carry_17_20));
wire w_sum_17_18, w_carry_17_18;
math_adder_full FA_17_18(.i_a(w_carry_16_20), .i_b(w_carry_16_18), .i_c(w_carry_16_16), .ow_sum(w_sum_17_18), .ow_carry(w_carry_17_18));
wire w_sum_17_16, w_carry_17_16;
math_adder_full FA_17_16(.i_a(w_carry_16_14), .i_b(w_carry_16_12), .i_c(w_carry_16_10), .ow_sum(w_sum_17_16), .ow_carry(w_carry_17_16));
wire w_sum_17_14, w_carry_17_14;
math_adder_full FA_17_14(.i_a(w_carry_16_08), .i_b(w_carry_16_06), .i_c(w_carry_16_04), .ow_sum(w_sum_17_14), .ow_carry(w_carry_17_14));
wire w_sum_17_12, w_carry_17_12;
math_adder_full FA_17_12(.i_a(w_carry_16_02), .i_b(w_sum_17_34), .i_c(w_sum_17_32), .ow_sum(w_sum_17_12), .ow_carry(w_carry_17_12));
wire w_sum_17_10, w_carry_17_10;
math_adder_full FA_17_10(.i_a(w_sum_17_30), .i_b(w_sum_17_28), .i_c(w_sum_17_26), .ow_sum(w_sum_17_10), .ow_carry(w_carry_17_10));
wire w_sum_17_08, w_carry_17_08;
math_adder_full FA_17_08(.i_a(w_sum_17_24), .i_b(w_sum_17_22), .i_c(w_sum_17_20), .ow_sum(w_sum_17_08), .ow_carry(w_carry_17_08));
wire w_sum_17_06, w_carry_17_06;
math_adder_full FA_17_06(.i_a(w_sum_17_18), .i_b(w_sum_17_16), .i_c(w_sum_17_14), .ow_sum(w_sum_17_06), .ow_carry(w_carry_17_06));
wire w_sum_17_04, w_carry_17_04;
math_adder_full FA_17_04(.i_a(w_sum_17_12), .i_b(w_sum_17_10), .i_c(w_sum_17_08), .ow_sum(w_sum_17_04), .ow_carry(w_carry_17_04));
wire w_sum_17_02, w_carry_17_02;
math_adder_half HA_17_02(.i_a(w_sum_17_06), .i_b(w_sum_17_04), .ow_sum(w_sum_17_02), .ow_carry(w_carry_17_02));
wire w_sum_18_36, w_carry_18_36;
math_adder_full FA_18_36(.i_a(w_pp_00_18), .i_b(w_pp_01_17), .i_c(w_pp_02_16), .ow_sum(w_sum_18_36), .ow_carry(w_carry_18_36));
wire w_sum_18_34, w_carry_18_34;
math_adder_full FA_18_34(.i_a(w_pp_03_15), .i_b(w_pp_04_14), .i_c(w_pp_05_13), .ow_sum(w_sum_18_34), .ow_carry(w_carry_18_34));
wire w_sum_18_32, w_carry_18_32;
math_adder_full FA_18_32(.i_a(w_pp_06_12), .i_b(w_pp_07_11), .i_c(w_pp_08_10), .ow_sum(w_sum_18_32), .ow_carry(w_carry_18_32));
wire w_sum_18_30, w_carry_18_30;
math_adder_full FA_18_30(.i_a(w_pp_09_09), .i_b(w_pp_10_08), .i_c(w_pp_11_07), .ow_sum(w_sum_18_30), .ow_carry(w_carry_18_30));
wire w_sum_18_28, w_carry_18_28;
math_adder_full FA_18_28(.i_a(w_pp_12_06), .i_b(w_pp_13_05), .i_c(w_pp_14_04), .ow_sum(w_sum_18_28), .ow_carry(w_carry_18_28));
wire w_sum_18_26, w_carry_18_26;
math_adder_full FA_18_26(.i_a(w_pp_15_03), .i_b(w_pp_16_02), .i_c(w_pp_17_01), .ow_sum(w_sum_18_26), .ow_carry(w_carry_18_26));
wire w_sum_18_24, w_carry_18_24;
math_adder_full FA_18_24(.i_a(w_pp_18_00), .i_b(w_carry_17_34), .i_c(w_carry_17_32), .ow_sum(w_sum_18_24), .ow_carry(w_carry_18_24));
wire w_sum_18_22, w_carry_18_22;
math_adder_full FA_18_22(.i_a(w_carry_17_30), .i_b(w_carry_17_28), .i_c(w_carry_17_26), .ow_sum(w_sum_18_22), .ow_carry(w_carry_18_22));
wire w_sum_18_20, w_carry_18_20;
math_adder_full FA_18_20(.i_a(w_carry_17_24), .i_b(w_carry_17_22), .i_c(w_carry_17_20), .ow_sum(w_sum_18_20), .ow_carry(w_carry_18_20));
wire w_sum_18_18, w_carry_18_18;
math_adder_full FA_18_18(.i_a(w_carry_17_18), .i_b(w_carry_17_16), .i_c(w_carry_17_14), .ow_sum(w_sum_18_18), .ow_carry(w_carry_18_18));
wire w_sum_18_16, w_carry_18_16;
math_adder_full FA_18_16(.i_a(w_carry_17_12), .i_b(w_carry_17_10), .i_c(w_carry_17_08), .ow_sum(w_sum_18_16), .ow_carry(w_carry_18_16));
wire w_sum_18_14, w_carry_18_14;
math_adder_full FA_18_14(.i_a(w_carry_17_06), .i_b(w_carry_17_04), .i_c(w_carry_17_02), .ow_sum(w_sum_18_14), .ow_carry(w_carry_18_14));
wire w_sum_18_12, w_carry_18_12;
math_adder_full FA_18_12(.i_a(w_sum_18_36), .i_b(w_sum_18_34), .i_c(w_sum_18_32), .ow_sum(w_sum_18_12), .ow_carry(w_carry_18_12));
wire w_sum_18_10, w_carry_18_10;
math_adder_full FA_18_10(.i_a(w_sum_18_30), .i_b(w_sum_18_28), .i_c(w_sum_18_26), .ow_sum(w_sum_18_10), .ow_carry(w_carry_18_10));
wire w_sum_18_08, w_carry_18_08;
math_adder_full FA_18_08(.i_a(w_sum_18_24), .i_b(w_sum_18_22), .i_c(w_sum_18_20), .ow_sum(w_sum_18_08), .ow_carry(w_carry_18_08));
wire w_sum_18_06, w_carry_18_06;
math_adder_full FA_18_06(.i_a(w_sum_18_18), .i_b(w_sum_18_16), .i_c(w_sum_18_14), .ow_sum(w_sum_18_06), .ow_carry(w_carry_18_06));
wire w_sum_18_04, w_carry_18_04;
math_adder_full FA_18_04(.i_a(w_sum_18_12), .i_b(w_sum_18_10), .i_c(w_sum_18_08), .ow_sum(w_sum_18_04), .ow_carry(w_carry_18_04));
wire w_sum_18_02, w_carry_18_02;
math_adder_half HA_18_02(.i_a(w_sum_18_06), .i_b(w_sum_18_04), .ow_sum(w_sum_18_02), .ow_carry(w_carry_18_02));
wire w_sum_19_38, w_carry_19_38;
math_adder_full FA_19_38(.i_a(w_pp_00_19), .i_b(w_pp_01_18), .i_c(w_pp_02_17), .ow_sum(w_sum_19_38), .ow_carry(w_carry_19_38));
wire w_sum_19_36, w_carry_19_36;
math_adder_full FA_19_36(.i_a(w_pp_03_16), .i_b(w_pp_04_15), .i_c(w_pp_05_14), .ow_sum(w_sum_19_36), .ow_carry(w_carry_19_36));
wire w_sum_19_34, w_carry_19_34;
math_adder_full FA_19_34(.i_a(w_pp_06_13), .i_b(w_pp_07_12), .i_c(w_pp_08_11), .ow_sum(w_sum_19_34), .ow_carry(w_carry_19_34));
wire w_sum_19_32, w_carry_19_32;
math_adder_full FA_19_32(.i_a(w_pp_09_10), .i_b(w_pp_10_09), .i_c(w_pp_11_08), .ow_sum(w_sum_19_32), .ow_carry(w_carry_19_32));
wire w_sum_19_30, w_carry_19_30;
math_adder_full FA_19_30(.i_a(w_pp_12_07), .i_b(w_pp_13_06), .i_c(w_pp_14_05), .ow_sum(w_sum_19_30), .ow_carry(w_carry_19_30));
wire w_sum_19_28, w_carry_19_28;
math_adder_full FA_19_28(.i_a(w_pp_15_04), .i_b(w_pp_16_03), .i_c(w_pp_17_02), .ow_sum(w_sum_19_28), .ow_carry(w_carry_19_28));
wire w_sum_19_26, w_carry_19_26;
math_adder_full FA_19_26(.i_a(w_pp_18_01), .i_b(w_pp_19_00), .i_c(w_carry_18_36), .ow_sum(w_sum_19_26), .ow_carry(w_carry_19_26));
wire w_sum_19_24, w_carry_19_24;
math_adder_full FA_19_24(.i_a(w_carry_18_34), .i_b(w_carry_18_32), .i_c(w_carry_18_30), .ow_sum(w_sum_19_24), .ow_carry(w_carry_19_24));
wire w_sum_19_22, w_carry_19_22;
math_adder_full FA_19_22(.i_a(w_carry_18_28), .i_b(w_carry_18_26), .i_c(w_carry_18_24), .ow_sum(w_sum_19_22), .ow_carry(w_carry_19_22));
wire w_sum_19_20, w_carry_19_20;
math_adder_full FA_19_20(.i_a(w_carry_18_22), .i_b(w_carry_18_20), .i_c(w_carry_18_18), .ow_sum(w_sum_19_20), .ow_carry(w_carry_19_20));
wire w_sum_19_18, w_carry_19_18;
math_adder_full FA_19_18(.i_a(w_carry_18_16), .i_b(w_carry_18_14), .i_c(w_carry_18_12), .ow_sum(w_sum_19_18), .ow_carry(w_carry_19_18));
wire w_sum_19_16, w_carry_19_16;
math_adder_full FA_19_16(.i_a(w_carry_18_10), .i_b(w_carry_18_08), .i_c(w_carry_18_06), .ow_sum(w_sum_19_16), .ow_carry(w_carry_19_16));
wire w_sum_19_14, w_carry_19_14;
math_adder_full FA_19_14(.i_a(w_carry_18_04), .i_b(w_carry_18_02), .i_c(w_sum_19_38), .ow_sum(w_sum_19_14), .ow_carry(w_carry_19_14));
wire w_sum_19_12, w_carry_19_12;
math_adder_full FA_19_12(.i_a(w_sum_19_36), .i_b(w_sum_19_34), .i_c(w_sum_19_32), .ow_sum(w_sum_19_12), .ow_carry(w_carry_19_12));
wire w_sum_19_10, w_carry_19_10;
math_adder_full FA_19_10(.i_a(w_sum_19_30), .i_b(w_sum_19_28), .i_c(w_sum_19_26), .ow_sum(w_sum_19_10), .ow_carry(w_carry_19_10));
wire w_sum_19_08, w_carry_19_08;
math_adder_full FA_19_08(.i_a(w_sum_19_24), .i_b(w_sum_19_22), .i_c(w_sum_19_20), .ow_sum(w_sum_19_08), .ow_carry(w_carry_19_08));
wire w_sum_19_06, w_carry_19_06;
math_adder_full FA_19_06(.i_a(w_sum_19_18), .i_b(w_sum_19_16), .i_c(w_sum_19_14), .ow_sum(w_sum_19_06), .ow_carry(w_carry_19_06));
wire w_sum_19_04, w_carry_19_04;
math_adder_full FA_19_04(.i_a(w_sum_19_12), .i_b(w_sum_19_10), .i_c(w_sum_19_08), .ow_sum(w_sum_19_04), .ow_carry(w_carry_19_04));
wire w_sum_19_02, w_carry_19_02;
math_adder_half HA_19_02(.i_a(w_sum_19_06), .i_b(w_sum_19_04), .ow_sum(w_sum_19_02), .ow_carry(w_carry_19_02));
wire w_sum_20_40, w_carry_20_40;
math_adder_full FA_20_40(.i_a(w_pp_00_20), .i_b(w_pp_01_19), .i_c(w_pp_02_18), .ow_sum(w_sum_20_40), .ow_carry(w_carry_20_40));
wire w_sum_20_38, w_carry_20_38;
math_adder_full FA_20_38(.i_a(w_pp_03_17), .i_b(w_pp_04_16), .i_c(w_pp_05_15), .ow_sum(w_sum_20_38), .ow_carry(w_carry_20_38));
wire w_sum_20_36, w_carry_20_36;
math_adder_full FA_20_36(.i_a(w_pp_06_14), .i_b(w_pp_07_13), .i_c(w_pp_08_12), .ow_sum(w_sum_20_36), .ow_carry(w_carry_20_36));
wire w_sum_20_34, w_carry_20_34;
math_adder_full FA_20_34(.i_a(w_pp_09_11), .i_b(w_pp_10_10), .i_c(w_pp_11_09), .ow_sum(w_sum_20_34), .ow_carry(w_carry_20_34));
wire w_sum_20_32, w_carry_20_32;
math_adder_full FA_20_32(.i_a(w_pp_12_08), .i_b(w_pp_13_07), .i_c(w_pp_14_06), .ow_sum(w_sum_20_32), .ow_carry(w_carry_20_32));
wire w_sum_20_30, w_carry_20_30;
math_adder_full FA_20_30(.i_a(w_pp_15_05), .i_b(w_pp_16_04), .i_c(w_pp_17_03), .ow_sum(w_sum_20_30), .ow_carry(w_carry_20_30));
wire w_sum_20_28, w_carry_20_28;
math_adder_full FA_20_28(.i_a(w_pp_18_02), .i_b(w_pp_19_01), .i_c(w_pp_20_00), .ow_sum(w_sum_20_28), .ow_carry(w_carry_20_28));
wire w_sum_20_26, w_carry_20_26;
math_adder_full FA_20_26(.i_a(w_carry_19_38), .i_b(w_carry_19_36), .i_c(w_carry_19_34), .ow_sum(w_sum_20_26), .ow_carry(w_carry_20_26));
wire w_sum_20_24, w_carry_20_24;
math_adder_full FA_20_24(.i_a(w_carry_19_32), .i_b(w_carry_19_30), .i_c(w_carry_19_28), .ow_sum(w_sum_20_24), .ow_carry(w_carry_20_24));
wire w_sum_20_22, w_carry_20_22;
math_adder_full FA_20_22(.i_a(w_carry_19_26), .i_b(w_carry_19_24), .i_c(w_carry_19_22), .ow_sum(w_sum_20_22), .ow_carry(w_carry_20_22));
wire w_sum_20_20, w_carry_20_20;
math_adder_full FA_20_20(.i_a(w_carry_19_20), .i_b(w_carry_19_18), .i_c(w_carry_19_16), .ow_sum(w_sum_20_20), .ow_carry(w_carry_20_20));
wire w_sum_20_18, w_carry_20_18;
math_adder_full FA_20_18(.i_a(w_carry_19_14), .i_b(w_carry_19_12), .i_c(w_carry_19_10), .ow_sum(w_sum_20_18), .ow_carry(w_carry_20_18));
wire w_sum_20_16, w_carry_20_16;
math_adder_full FA_20_16(.i_a(w_carry_19_08), .i_b(w_carry_19_06), .i_c(w_carry_19_04), .ow_sum(w_sum_20_16), .ow_carry(w_carry_20_16));
wire w_sum_20_14, w_carry_20_14;
math_adder_full FA_20_14(.i_a(w_carry_19_02), .i_b(w_sum_20_40), .i_c(w_sum_20_38), .ow_sum(w_sum_20_14), .ow_carry(w_carry_20_14));
wire w_sum_20_12, w_carry_20_12;
math_adder_full FA_20_12(.i_a(w_sum_20_36), .i_b(w_sum_20_34), .i_c(w_sum_20_32), .ow_sum(w_sum_20_12), .ow_carry(w_carry_20_12));
wire w_sum_20_10, w_carry_20_10;
math_adder_full FA_20_10(.i_a(w_sum_20_30), .i_b(w_sum_20_28), .i_c(w_sum_20_26), .ow_sum(w_sum_20_10), .ow_carry(w_carry_20_10));
wire w_sum_20_08, w_carry_20_08;
math_adder_full FA_20_08(.i_a(w_sum_20_24), .i_b(w_sum_20_22), .i_c(w_sum_20_20), .ow_sum(w_sum_20_08), .ow_carry(w_carry_20_08));
wire w_sum_20_06, w_carry_20_06;
math_adder_full FA_20_06(.i_a(w_sum_20_18), .i_b(w_sum_20_16), .i_c(w_sum_20_14), .ow_sum(w_sum_20_06), .ow_carry(w_carry_20_06));
wire w_sum_20_04, w_carry_20_04;
math_adder_full FA_20_04(.i_a(w_sum_20_12), .i_b(w_sum_20_10), .i_c(w_sum_20_08), .ow_sum(w_sum_20_04), .ow_carry(w_carry_20_04));
wire w_sum_20_02, w_carry_20_02;
math_adder_half HA_20_02(.i_a(w_sum_20_06), .i_b(w_sum_20_04), .ow_sum(w_sum_20_02), .ow_carry(w_carry_20_02));
wire w_sum_21_42, w_carry_21_42;
math_adder_full FA_21_42(.i_a(w_pp_00_21), .i_b(w_pp_01_20), .i_c(w_pp_02_19), .ow_sum(w_sum_21_42), .ow_carry(w_carry_21_42));
wire w_sum_21_40, w_carry_21_40;
math_adder_full FA_21_40(.i_a(w_pp_03_18), .i_b(w_pp_04_17), .i_c(w_pp_05_16), .ow_sum(w_sum_21_40), .ow_carry(w_carry_21_40));
wire w_sum_21_38, w_carry_21_38;
math_adder_full FA_21_38(.i_a(w_pp_06_15), .i_b(w_pp_07_14), .i_c(w_pp_08_13), .ow_sum(w_sum_21_38), .ow_carry(w_carry_21_38));
wire w_sum_21_36, w_carry_21_36;
math_adder_full FA_21_36(.i_a(w_pp_09_12), .i_b(w_pp_10_11), .i_c(w_pp_11_10), .ow_sum(w_sum_21_36), .ow_carry(w_carry_21_36));
wire w_sum_21_34, w_carry_21_34;
math_adder_full FA_21_34(.i_a(w_pp_12_09), .i_b(w_pp_13_08), .i_c(w_pp_14_07), .ow_sum(w_sum_21_34), .ow_carry(w_carry_21_34));
wire w_sum_21_32, w_carry_21_32;
math_adder_full FA_21_32(.i_a(w_pp_15_06), .i_b(w_pp_16_05), .i_c(w_pp_17_04), .ow_sum(w_sum_21_32), .ow_carry(w_carry_21_32));
wire w_sum_21_30, w_carry_21_30;
math_adder_full FA_21_30(.i_a(w_pp_18_03), .i_b(w_pp_19_02), .i_c(w_pp_20_01), .ow_sum(w_sum_21_30), .ow_carry(w_carry_21_30));
wire w_sum_21_28, w_carry_21_28;
math_adder_full FA_21_28(.i_a(w_pp_21_00), .i_b(w_carry_20_40), .i_c(w_carry_20_38), .ow_sum(w_sum_21_28), .ow_carry(w_carry_21_28));
wire w_sum_21_26, w_carry_21_26;
math_adder_full FA_21_26(.i_a(w_carry_20_36), .i_b(w_carry_20_34), .i_c(w_carry_20_32), .ow_sum(w_sum_21_26), .ow_carry(w_carry_21_26));
wire w_sum_21_24, w_carry_21_24;
math_adder_full FA_21_24(.i_a(w_carry_20_30), .i_b(w_carry_20_28), .i_c(w_carry_20_26), .ow_sum(w_sum_21_24), .ow_carry(w_carry_21_24));
wire w_sum_21_22, w_carry_21_22;
math_adder_full FA_21_22(.i_a(w_carry_20_24), .i_b(w_carry_20_22), .i_c(w_carry_20_20), .ow_sum(w_sum_21_22), .ow_carry(w_carry_21_22));
wire w_sum_21_20, w_carry_21_20;
math_adder_full FA_21_20(.i_a(w_carry_20_18), .i_b(w_carry_20_16), .i_c(w_carry_20_14), .ow_sum(w_sum_21_20), .ow_carry(w_carry_21_20));
wire w_sum_21_18, w_carry_21_18;
math_adder_full FA_21_18(.i_a(w_carry_20_12), .i_b(w_carry_20_10), .i_c(w_carry_20_08), .ow_sum(w_sum_21_18), .ow_carry(w_carry_21_18));
wire w_sum_21_16, w_carry_21_16;
math_adder_full FA_21_16(.i_a(w_carry_20_06), .i_b(w_carry_20_04), .i_c(w_carry_20_02), .ow_sum(w_sum_21_16), .ow_carry(w_carry_21_16));
wire w_sum_21_14, w_carry_21_14;
math_adder_full FA_21_14(.i_a(w_sum_21_42), .i_b(w_sum_21_40), .i_c(w_sum_21_38), .ow_sum(w_sum_21_14), .ow_carry(w_carry_21_14));
wire w_sum_21_12, w_carry_21_12;
math_adder_full FA_21_12(.i_a(w_sum_21_36), .i_b(w_sum_21_34), .i_c(w_sum_21_32), .ow_sum(w_sum_21_12), .ow_carry(w_carry_21_12));
wire w_sum_21_10, w_carry_21_10;
math_adder_full FA_21_10(.i_a(w_sum_21_30), .i_b(w_sum_21_28), .i_c(w_sum_21_26), .ow_sum(w_sum_21_10), .ow_carry(w_carry_21_10));
wire w_sum_21_08, w_carry_21_08;
math_adder_full FA_21_08(.i_a(w_sum_21_24), .i_b(w_sum_21_22), .i_c(w_sum_21_20), .ow_sum(w_sum_21_08), .ow_carry(w_carry_21_08));
wire w_sum_21_06, w_carry_21_06;
math_adder_full FA_21_06(.i_a(w_sum_21_18), .i_b(w_sum_21_16), .i_c(w_sum_21_14), .ow_sum(w_sum_21_06), .ow_carry(w_carry_21_06));
wire w_sum_21_04, w_carry_21_04;
math_adder_full FA_21_04(.i_a(w_sum_21_12), .i_b(w_sum_21_10), .i_c(w_sum_21_08), .ow_sum(w_sum_21_04), .ow_carry(w_carry_21_04));
wire w_sum_21_02, w_carry_21_02;
math_adder_half HA_21_02(.i_a(w_sum_21_06), .i_b(w_sum_21_04), .ow_sum(w_sum_21_02), .ow_carry(w_carry_21_02));
wire w_sum_22_44, w_carry_22_44;
math_adder_full FA_22_44(.i_a(w_pp_00_22), .i_b(w_pp_01_21), .i_c(w_pp_02_20), .ow_sum(w_sum_22_44), .ow_carry(w_carry_22_44));
wire w_sum_22_42, w_carry_22_42;
math_adder_full FA_22_42(.i_a(w_pp_03_19), .i_b(w_pp_04_18), .i_c(w_pp_05_17), .ow_sum(w_sum_22_42), .ow_carry(w_carry_22_42));
wire w_sum_22_40, w_carry_22_40;
math_adder_full FA_22_40(.i_a(w_pp_06_16), .i_b(w_pp_07_15), .i_c(w_pp_08_14), .ow_sum(w_sum_22_40), .ow_carry(w_carry_22_40));
wire w_sum_22_38, w_carry_22_38;
math_adder_full FA_22_38(.i_a(w_pp_09_13), .i_b(w_pp_10_12), .i_c(w_pp_11_11), .ow_sum(w_sum_22_38), .ow_carry(w_carry_22_38));
wire w_sum_22_36, w_carry_22_36;
math_adder_full FA_22_36(.i_a(w_pp_12_10), .i_b(w_pp_13_09), .i_c(w_pp_14_08), .ow_sum(w_sum_22_36), .ow_carry(w_carry_22_36));
wire w_sum_22_34, w_carry_22_34;
math_adder_full FA_22_34(.i_a(w_pp_15_07), .i_b(w_pp_16_06), .i_c(w_pp_17_05), .ow_sum(w_sum_22_34), .ow_carry(w_carry_22_34));
wire w_sum_22_32, w_carry_22_32;
math_adder_full FA_22_32(.i_a(w_pp_18_04), .i_b(w_pp_19_03), .i_c(w_pp_20_02), .ow_sum(w_sum_22_32), .ow_carry(w_carry_22_32));
wire w_sum_22_30, w_carry_22_30;
math_adder_full FA_22_30(.i_a(w_pp_21_01), .i_b(w_pp_22_00), .i_c(w_carry_21_42), .ow_sum(w_sum_22_30), .ow_carry(w_carry_22_30));
wire w_sum_22_28, w_carry_22_28;
math_adder_full FA_22_28(.i_a(w_carry_21_40), .i_b(w_carry_21_38), .i_c(w_carry_21_36), .ow_sum(w_sum_22_28), .ow_carry(w_carry_22_28));
wire w_sum_22_26, w_carry_22_26;
math_adder_full FA_22_26(.i_a(w_carry_21_34), .i_b(w_carry_21_32), .i_c(w_carry_21_30), .ow_sum(w_sum_22_26), .ow_carry(w_carry_22_26));
wire w_sum_22_24, w_carry_22_24;
math_adder_full FA_22_24(.i_a(w_carry_21_28), .i_b(w_carry_21_26), .i_c(w_carry_21_24), .ow_sum(w_sum_22_24), .ow_carry(w_carry_22_24));
wire w_sum_22_22, w_carry_22_22;
math_adder_full FA_22_22(.i_a(w_carry_21_22), .i_b(w_carry_21_20), .i_c(w_carry_21_18), .ow_sum(w_sum_22_22), .ow_carry(w_carry_22_22));
wire w_sum_22_20, w_carry_22_20;
math_adder_full FA_22_20(.i_a(w_carry_21_16), .i_b(w_carry_21_14), .i_c(w_carry_21_12), .ow_sum(w_sum_22_20), .ow_carry(w_carry_22_20));
wire w_sum_22_18, w_carry_22_18;
math_adder_full FA_22_18(.i_a(w_carry_21_10), .i_b(w_carry_21_08), .i_c(w_carry_21_06), .ow_sum(w_sum_22_18), .ow_carry(w_carry_22_18));
wire w_sum_22_16, w_carry_22_16;
math_adder_full FA_22_16(.i_a(w_carry_21_04), .i_b(w_carry_21_02), .i_c(w_sum_22_44), .ow_sum(w_sum_22_16), .ow_carry(w_carry_22_16));
wire w_sum_22_14, w_carry_22_14;
math_adder_full FA_22_14(.i_a(w_sum_22_42), .i_b(w_sum_22_40), .i_c(w_sum_22_38), .ow_sum(w_sum_22_14), .ow_carry(w_carry_22_14));
wire w_sum_22_12, w_carry_22_12;
math_adder_full FA_22_12(.i_a(w_sum_22_36), .i_b(w_sum_22_34), .i_c(w_sum_22_32), .ow_sum(w_sum_22_12), .ow_carry(w_carry_22_12));
wire w_sum_22_10, w_carry_22_10;
math_adder_full FA_22_10(.i_a(w_sum_22_30), .i_b(w_sum_22_28), .i_c(w_sum_22_26), .ow_sum(w_sum_22_10), .ow_carry(w_carry_22_10));
wire w_sum_22_08, w_carry_22_08;
math_adder_full FA_22_08(.i_a(w_sum_22_24), .i_b(w_sum_22_22), .i_c(w_sum_22_20), .ow_sum(w_sum_22_08), .ow_carry(w_carry_22_08));
wire w_sum_22_06, w_carry_22_06;
math_adder_full FA_22_06(.i_a(w_sum_22_18), .i_b(w_sum_22_16), .i_c(w_sum_22_14), .ow_sum(w_sum_22_06), .ow_carry(w_carry_22_06));
wire w_sum_22_04, w_carry_22_04;
math_adder_full FA_22_04(.i_a(w_sum_22_12), .i_b(w_sum_22_10), .i_c(w_sum_22_08), .ow_sum(w_sum_22_04), .ow_carry(w_carry_22_04));
wire w_sum_22_02, w_carry_22_02;
math_adder_half HA_22_02(.i_a(w_sum_22_06), .i_b(w_sum_22_04), .ow_sum(w_sum_22_02), .ow_carry(w_carry_22_02));
wire w_sum_23_46, w_carry_23_46;
math_adder_full FA_23_46(.i_a(w_pp_00_23), .i_b(w_pp_01_22), .i_c(w_pp_02_21), .ow_sum(w_sum_23_46), .ow_carry(w_carry_23_46));
wire w_sum_23_44, w_carry_23_44;
math_adder_full FA_23_44(.i_a(w_pp_03_20), .i_b(w_pp_04_19), .i_c(w_pp_05_18), .ow_sum(w_sum_23_44), .ow_carry(w_carry_23_44));
wire w_sum_23_42, w_carry_23_42;
math_adder_full FA_23_42(.i_a(w_pp_06_17), .i_b(w_pp_07_16), .i_c(w_pp_08_15), .ow_sum(w_sum_23_42), .ow_carry(w_carry_23_42));
wire w_sum_23_40, w_carry_23_40;
math_adder_full FA_23_40(.i_a(w_pp_09_14), .i_b(w_pp_10_13), .i_c(w_pp_11_12), .ow_sum(w_sum_23_40), .ow_carry(w_carry_23_40));
wire w_sum_23_38, w_carry_23_38;
math_adder_full FA_23_38(.i_a(w_pp_12_11), .i_b(w_pp_13_10), .i_c(w_pp_14_09), .ow_sum(w_sum_23_38), .ow_carry(w_carry_23_38));
wire w_sum_23_36, w_carry_23_36;
math_adder_full FA_23_36(.i_a(w_pp_15_08), .i_b(w_pp_16_07), .i_c(w_pp_17_06), .ow_sum(w_sum_23_36), .ow_carry(w_carry_23_36));
wire w_sum_23_34, w_carry_23_34;
math_adder_full FA_23_34(.i_a(w_pp_18_05), .i_b(w_pp_19_04), .i_c(w_pp_20_03), .ow_sum(w_sum_23_34), .ow_carry(w_carry_23_34));
wire w_sum_23_32, w_carry_23_32;
math_adder_full FA_23_32(.i_a(w_pp_21_02), .i_b(w_pp_22_01), .i_c(w_pp_23_00), .ow_sum(w_sum_23_32), .ow_carry(w_carry_23_32));
wire w_sum_23_30, w_carry_23_30;
math_adder_full FA_23_30(.i_a(w_carry_22_44), .i_b(w_carry_22_42), .i_c(w_carry_22_40), .ow_sum(w_sum_23_30), .ow_carry(w_carry_23_30));
wire w_sum_23_28, w_carry_23_28;
math_adder_full FA_23_28(.i_a(w_carry_22_38), .i_b(w_carry_22_36), .i_c(w_carry_22_34), .ow_sum(w_sum_23_28), .ow_carry(w_carry_23_28));
wire w_sum_23_26, w_carry_23_26;
math_adder_full FA_23_26(.i_a(w_carry_22_32), .i_b(w_carry_22_30), .i_c(w_carry_22_28), .ow_sum(w_sum_23_26), .ow_carry(w_carry_23_26));
wire w_sum_23_24, w_carry_23_24;
math_adder_full FA_23_24(.i_a(w_carry_22_26), .i_b(w_carry_22_24), .i_c(w_carry_22_22), .ow_sum(w_sum_23_24), .ow_carry(w_carry_23_24));
wire w_sum_23_22, w_carry_23_22;
math_adder_full FA_23_22(.i_a(w_carry_22_20), .i_b(w_carry_22_18), .i_c(w_carry_22_16), .ow_sum(w_sum_23_22), .ow_carry(w_carry_23_22));
wire w_sum_23_20, w_carry_23_20;
math_adder_full FA_23_20(.i_a(w_carry_22_14), .i_b(w_carry_22_12), .i_c(w_carry_22_10), .ow_sum(w_sum_23_20), .ow_carry(w_carry_23_20));
wire w_sum_23_18, w_carry_23_18;
math_adder_full FA_23_18(.i_a(w_carry_22_08), .i_b(w_carry_22_06), .i_c(w_carry_22_04), .ow_sum(w_sum_23_18), .ow_carry(w_carry_23_18));
wire w_sum_23_16, w_carry_23_16;
math_adder_full FA_23_16(.i_a(w_carry_22_02), .i_b(w_sum_23_46), .i_c(w_sum_23_44), .ow_sum(w_sum_23_16), .ow_carry(w_carry_23_16));
wire w_sum_23_14, w_carry_23_14;
math_adder_full FA_23_14(.i_a(w_sum_23_42), .i_b(w_sum_23_40), .i_c(w_sum_23_38), .ow_sum(w_sum_23_14), .ow_carry(w_carry_23_14));
wire w_sum_23_12, w_carry_23_12;
math_adder_full FA_23_12(.i_a(w_sum_23_36), .i_b(w_sum_23_34), .i_c(w_sum_23_32), .ow_sum(w_sum_23_12), .ow_carry(w_carry_23_12));
wire w_sum_23_10, w_carry_23_10;
math_adder_full FA_23_10(.i_a(w_sum_23_30), .i_b(w_sum_23_28), .i_c(w_sum_23_26), .ow_sum(w_sum_23_10), .ow_carry(w_carry_23_10));
wire w_sum_23_08, w_carry_23_08;
math_adder_full FA_23_08(.i_a(w_sum_23_24), .i_b(w_sum_23_22), .i_c(w_sum_23_20), .ow_sum(w_sum_23_08), .ow_carry(w_carry_23_08));
wire w_sum_23_06, w_carry_23_06;
math_adder_full FA_23_06(.i_a(w_sum_23_18), .i_b(w_sum_23_16), .i_c(w_sum_23_14), .ow_sum(w_sum_23_06), .ow_carry(w_carry_23_06));
wire w_sum_23_04, w_carry_23_04;
math_adder_full FA_23_04(.i_a(w_sum_23_12), .i_b(w_sum_23_10), .i_c(w_sum_23_08), .ow_sum(w_sum_23_04), .ow_carry(w_carry_23_04));
wire w_sum_23_02, w_carry_23_02;
math_adder_half HA_23_02(.i_a(w_sum_23_06), .i_b(w_sum_23_04), .ow_sum(w_sum_23_02), .ow_carry(w_carry_23_02));
wire w_sum_24_48, w_carry_24_48;
math_adder_full FA_24_48(.i_a(w_pp_00_24), .i_b(w_pp_01_23), .i_c(w_pp_02_22), .ow_sum(w_sum_24_48), .ow_carry(w_carry_24_48));
wire w_sum_24_46, w_carry_24_46;
math_adder_full FA_24_46(.i_a(w_pp_03_21), .i_b(w_pp_04_20), .i_c(w_pp_05_19), .ow_sum(w_sum_24_46), .ow_carry(w_carry_24_46));
wire w_sum_24_44, w_carry_24_44;
math_adder_full FA_24_44(.i_a(w_pp_06_18), .i_b(w_pp_07_17), .i_c(w_pp_08_16), .ow_sum(w_sum_24_44), .ow_carry(w_carry_24_44));
wire w_sum_24_42, w_carry_24_42;
math_adder_full FA_24_42(.i_a(w_pp_09_15), .i_b(w_pp_10_14), .i_c(w_pp_11_13), .ow_sum(w_sum_24_42), .ow_carry(w_carry_24_42));
wire w_sum_24_40, w_carry_24_40;
math_adder_full FA_24_40(.i_a(w_pp_12_12), .i_b(w_pp_13_11), .i_c(w_pp_14_10), .ow_sum(w_sum_24_40), .ow_carry(w_carry_24_40));
wire w_sum_24_38, w_carry_24_38;
math_adder_full FA_24_38(.i_a(w_pp_15_09), .i_b(w_pp_16_08), .i_c(w_pp_17_07), .ow_sum(w_sum_24_38), .ow_carry(w_carry_24_38));
wire w_sum_24_36, w_carry_24_36;
math_adder_full FA_24_36(.i_a(w_pp_18_06), .i_b(w_pp_19_05), .i_c(w_pp_20_04), .ow_sum(w_sum_24_36), .ow_carry(w_carry_24_36));
wire w_sum_24_34, w_carry_24_34;
math_adder_full FA_24_34(.i_a(w_pp_21_03), .i_b(w_pp_22_02), .i_c(w_pp_23_01), .ow_sum(w_sum_24_34), .ow_carry(w_carry_24_34));
wire w_sum_24_32, w_carry_24_32;
math_adder_full FA_24_32(.i_a(w_pp_24_00), .i_b(w_carry_23_46), .i_c(w_carry_23_44), .ow_sum(w_sum_24_32), .ow_carry(w_carry_24_32));
wire w_sum_24_30, w_carry_24_30;
math_adder_full FA_24_30(.i_a(w_carry_23_42), .i_b(w_carry_23_40), .i_c(w_carry_23_38), .ow_sum(w_sum_24_30), .ow_carry(w_carry_24_30));
wire w_sum_24_28, w_carry_24_28;
math_adder_full FA_24_28(.i_a(w_carry_23_36), .i_b(w_carry_23_34), .i_c(w_carry_23_32), .ow_sum(w_sum_24_28), .ow_carry(w_carry_24_28));
wire w_sum_24_26, w_carry_24_26;
math_adder_full FA_24_26(.i_a(w_carry_23_30), .i_b(w_carry_23_28), .i_c(w_carry_23_26), .ow_sum(w_sum_24_26), .ow_carry(w_carry_24_26));
wire w_sum_24_24, w_carry_24_24;
math_adder_full FA_24_24(.i_a(w_carry_23_24), .i_b(w_carry_23_22), .i_c(w_carry_23_20), .ow_sum(w_sum_24_24), .ow_carry(w_carry_24_24));
wire w_sum_24_22, w_carry_24_22;
math_adder_full FA_24_22(.i_a(w_carry_23_18), .i_b(w_carry_23_16), .i_c(w_carry_23_14), .ow_sum(w_sum_24_22), .ow_carry(w_carry_24_22));
wire w_sum_24_20, w_carry_24_20;
math_adder_full FA_24_20(.i_a(w_carry_23_12), .i_b(w_carry_23_10), .i_c(w_carry_23_08), .ow_sum(w_sum_24_20), .ow_carry(w_carry_24_20));
wire w_sum_24_18, w_carry_24_18;
math_adder_full FA_24_18(.i_a(w_carry_23_06), .i_b(w_carry_23_04), .i_c(w_carry_23_02), .ow_sum(w_sum_24_18), .ow_carry(w_carry_24_18));
wire w_sum_24_16, w_carry_24_16;
math_adder_full FA_24_16(.i_a(w_sum_24_48), .i_b(w_sum_24_46), .i_c(w_sum_24_44), .ow_sum(w_sum_24_16), .ow_carry(w_carry_24_16));
wire w_sum_24_14, w_carry_24_14;
math_adder_full FA_24_14(.i_a(w_sum_24_42), .i_b(w_sum_24_40), .i_c(w_sum_24_38), .ow_sum(w_sum_24_14), .ow_carry(w_carry_24_14));
wire w_sum_24_12, w_carry_24_12;
math_adder_full FA_24_12(.i_a(w_sum_24_36), .i_b(w_sum_24_34), .i_c(w_sum_24_32), .ow_sum(w_sum_24_12), .ow_carry(w_carry_24_12));
wire w_sum_24_10, w_carry_24_10;
math_adder_full FA_24_10(.i_a(w_sum_24_30), .i_b(w_sum_24_28), .i_c(w_sum_24_26), .ow_sum(w_sum_24_10), .ow_carry(w_carry_24_10));
wire w_sum_24_08, w_carry_24_08;
math_adder_full FA_24_08(.i_a(w_sum_24_24), .i_b(w_sum_24_22), .i_c(w_sum_24_20), .ow_sum(w_sum_24_08), .ow_carry(w_carry_24_08));
wire w_sum_24_06, w_carry_24_06;
math_adder_full FA_24_06(.i_a(w_sum_24_18), .i_b(w_sum_24_16), .i_c(w_sum_24_14), .ow_sum(w_sum_24_06), .ow_carry(w_carry_24_06));
wire w_sum_24_04, w_carry_24_04;
math_adder_full FA_24_04(.i_a(w_sum_24_12), .i_b(w_sum_24_10), .i_c(w_sum_24_08), .ow_sum(w_sum_24_04), .ow_carry(w_carry_24_04));
wire w_sum_24_02, w_carry_24_02;
math_adder_half HA_24_02(.i_a(w_sum_24_06), .i_b(w_sum_24_04), .ow_sum(w_sum_24_02), .ow_carry(w_carry_24_02));
wire w_sum_25_50, w_carry_25_50;
math_adder_full FA_25_50(.i_a(w_pp_00_25), .i_b(w_pp_01_24), .i_c(w_pp_02_23), .ow_sum(w_sum_25_50), .ow_carry(w_carry_25_50));
wire w_sum_25_48, w_carry_25_48;
math_adder_full FA_25_48(.i_a(w_pp_03_22), .i_b(w_pp_04_21), .i_c(w_pp_05_20), .ow_sum(w_sum_25_48), .ow_carry(w_carry_25_48));
wire w_sum_25_46, w_carry_25_46;
math_adder_full FA_25_46(.i_a(w_pp_06_19), .i_b(w_pp_07_18), .i_c(w_pp_08_17), .ow_sum(w_sum_25_46), .ow_carry(w_carry_25_46));
wire w_sum_25_44, w_carry_25_44;
math_adder_full FA_25_44(.i_a(w_pp_09_16), .i_b(w_pp_10_15), .i_c(w_pp_11_14), .ow_sum(w_sum_25_44), .ow_carry(w_carry_25_44));
wire w_sum_25_42, w_carry_25_42;
math_adder_full FA_25_42(.i_a(w_pp_12_13), .i_b(w_pp_13_12), .i_c(w_pp_14_11), .ow_sum(w_sum_25_42), .ow_carry(w_carry_25_42));
wire w_sum_25_40, w_carry_25_40;
math_adder_full FA_25_40(.i_a(w_pp_15_10), .i_b(w_pp_16_09), .i_c(w_pp_17_08), .ow_sum(w_sum_25_40), .ow_carry(w_carry_25_40));
wire w_sum_25_38, w_carry_25_38;
math_adder_full FA_25_38(.i_a(w_pp_18_07), .i_b(w_pp_19_06), .i_c(w_pp_20_05), .ow_sum(w_sum_25_38), .ow_carry(w_carry_25_38));
wire w_sum_25_36, w_carry_25_36;
math_adder_full FA_25_36(.i_a(w_pp_21_04), .i_b(w_pp_22_03), .i_c(w_pp_23_02), .ow_sum(w_sum_25_36), .ow_carry(w_carry_25_36));
wire w_sum_25_34, w_carry_25_34;
math_adder_full FA_25_34(.i_a(w_pp_24_01), .i_b(w_pp_25_00), .i_c(w_carry_24_48), .ow_sum(w_sum_25_34), .ow_carry(w_carry_25_34));
wire w_sum_25_32, w_carry_25_32;
math_adder_full FA_25_32(.i_a(w_carry_24_46), .i_b(w_carry_24_44), .i_c(w_carry_24_42), .ow_sum(w_sum_25_32), .ow_carry(w_carry_25_32));
wire w_sum_25_30, w_carry_25_30;
math_adder_full FA_25_30(.i_a(w_carry_24_40), .i_b(w_carry_24_38), .i_c(w_carry_24_36), .ow_sum(w_sum_25_30), .ow_carry(w_carry_25_30));
wire w_sum_25_28, w_carry_25_28;
math_adder_full FA_25_28(.i_a(w_carry_24_34), .i_b(w_carry_24_32), .i_c(w_carry_24_30), .ow_sum(w_sum_25_28), .ow_carry(w_carry_25_28));
wire w_sum_25_26, w_carry_25_26;
math_adder_full FA_25_26(.i_a(w_carry_24_28), .i_b(w_carry_24_26), .i_c(w_carry_24_24), .ow_sum(w_sum_25_26), .ow_carry(w_carry_25_26));
wire w_sum_25_24, w_carry_25_24;
math_adder_full FA_25_24(.i_a(w_carry_24_22), .i_b(w_carry_24_20), .i_c(w_carry_24_18), .ow_sum(w_sum_25_24), .ow_carry(w_carry_25_24));
wire w_sum_25_22, w_carry_25_22;
math_adder_full FA_25_22(.i_a(w_carry_24_16), .i_b(w_carry_24_14), .i_c(w_carry_24_12), .ow_sum(w_sum_25_22), .ow_carry(w_carry_25_22));
wire w_sum_25_20, w_carry_25_20;
math_adder_full FA_25_20(.i_a(w_carry_24_10), .i_b(w_carry_24_08), .i_c(w_carry_24_06), .ow_sum(w_sum_25_20), .ow_carry(w_carry_25_20));
wire w_sum_25_18, w_carry_25_18;
math_adder_full FA_25_18(.i_a(w_carry_24_04), .i_b(w_carry_24_02), .i_c(w_sum_25_50), .ow_sum(w_sum_25_18), .ow_carry(w_carry_25_18));
wire w_sum_25_16, w_carry_25_16;
math_adder_full FA_25_16(.i_a(w_sum_25_48), .i_b(w_sum_25_46), .i_c(w_sum_25_44), .ow_sum(w_sum_25_16), .ow_carry(w_carry_25_16));
wire w_sum_25_14, w_carry_25_14;
math_adder_full FA_25_14(.i_a(w_sum_25_42), .i_b(w_sum_25_40), .i_c(w_sum_25_38), .ow_sum(w_sum_25_14), .ow_carry(w_carry_25_14));
wire w_sum_25_12, w_carry_25_12;
math_adder_full FA_25_12(.i_a(w_sum_25_36), .i_b(w_sum_25_34), .i_c(w_sum_25_32), .ow_sum(w_sum_25_12), .ow_carry(w_carry_25_12));
wire w_sum_25_10, w_carry_25_10;
math_adder_full FA_25_10(.i_a(w_sum_25_30), .i_b(w_sum_25_28), .i_c(w_sum_25_26), .ow_sum(w_sum_25_10), .ow_carry(w_carry_25_10));
wire w_sum_25_08, w_carry_25_08;
math_adder_full FA_25_08(.i_a(w_sum_25_24), .i_b(w_sum_25_22), .i_c(w_sum_25_20), .ow_sum(w_sum_25_08), .ow_carry(w_carry_25_08));
wire w_sum_25_06, w_carry_25_06;
math_adder_full FA_25_06(.i_a(w_sum_25_18), .i_b(w_sum_25_16), .i_c(w_sum_25_14), .ow_sum(w_sum_25_06), .ow_carry(w_carry_25_06));
wire w_sum_25_04, w_carry_25_04;
math_adder_full FA_25_04(.i_a(w_sum_25_12), .i_b(w_sum_25_10), .i_c(w_sum_25_08), .ow_sum(w_sum_25_04), .ow_carry(w_carry_25_04));
wire w_sum_25_02, w_carry_25_02;
math_adder_half HA_25_02(.i_a(w_sum_25_06), .i_b(w_sum_25_04), .ow_sum(w_sum_25_02), .ow_carry(w_carry_25_02));
wire w_sum_26_52, w_carry_26_52;
math_adder_full FA_26_52(.i_a(w_pp_00_26), .i_b(w_pp_01_25), .i_c(w_pp_02_24), .ow_sum(w_sum_26_52), .ow_carry(w_carry_26_52));
wire w_sum_26_50, w_carry_26_50;
math_adder_full FA_26_50(.i_a(w_pp_03_23), .i_b(w_pp_04_22), .i_c(w_pp_05_21), .ow_sum(w_sum_26_50), .ow_carry(w_carry_26_50));
wire w_sum_26_48, w_carry_26_48;
math_adder_full FA_26_48(.i_a(w_pp_06_20), .i_b(w_pp_07_19), .i_c(w_pp_08_18), .ow_sum(w_sum_26_48), .ow_carry(w_carry_26_48));
wire w_sum_26_46, w_carry_26_46;
math_adder_full FA_26_46(.i_a(w_pp_09_17), .i_b(w_pp_10_16), .i_c(w_pp_11_15), .ow_sum(w_sum_26_46), .ow_carry(w_carry_26_46));
wire w_sum_26_44, w_carry_26_44;
math_adder_full FA_26_44(.i_a(w_pp_12_14), .i_b(w_pp_13_13), .i_c(w_pp_14_12), .ow_sum(w_sum_26_44), .ow_carry(w_carry_26_44));
wire w_sum_26_42, w_carry_26_42;
math_adder_full FA_26_42(.i_a(w_pp_15_11), .i_b(w_pp_16_10), .i_c(w_pp_17_09), .ow_sum(w_sum_26_42), .ow_carry(w_carry_26_42));
wire w_sum_26_40, w_carry_26_40;
math_adder_full FA_26_40(.i_a(w_pp_18_08), .i_b(w_pp_19_07), .i_c(w_pp_20_06), .ow_sum(w_sum_26_40), .ow_carry(w_carry_26_40));
wire w_sum_26_38, w_carry_26_38;
math_adder_full FA_26_38(.i_a(w_pp_21_05), .i_b(w_pp_22_04), .i_c(w_pp_23_03), .ow_sum(w_sum_26_38), .ow_carry(w_carry_26_38));
wire w_sum_26_36, w_carry_26_36;
math_adder_full FA_26_36(.i_a(w_pp_24_02), .i_b(w_pp_25_01), .i_c(w_pp_26_00), .ow_sum(w_sum_26_36), .ow_carry(w_carry_26_36));
wire w_sum_26_34, w_carry_26_34;
math_adder_full FA_26_34(.i_a(w_carry_25_50), .i_b(w_carry_25_48), .i_c(w_carry_25_46), .ow_sum(w_sum_26_34), .ow_carry(w_carry_26_34));
wire w_sum_26_32, w_carry_26_32;
math_adder_full FA_26_32(.i_a(w_carry_25_44), .i_b(w_carry_25_42), .i_c(w_carry_25_40), .ow_sum(w_sum_26_32), .ow_carry(w_carry_26_32));
wire w_sum_26_30, w_carry_26_30;
math_adder_full FA_26_30(.i_a(w_carry_25_38), .i_b(w_carry_25_36), .i_c(w_carry_25_34), .ow_sum(w_sum_26_30), .ow_carry(w_carry_26_30));
wire w_sum_26_28, w_carry_26_28;
math_adder_full FA_26_28(.i_a(w_carry_25_32), .i_b(w_carry_25_30), .i_c(w_carry_25_28), .ow_sum(w_sum_26_28), .ow_carry(w_carry_26_28));
wire w_sum_26_26, w_carry_26_26;
math_adder_full FA_26_26(.i_a(w_carry_25_26), .i_b(w_carry_25_24), .i_c(w_carry_25_22), .ow_sum(w_sum_26_26), .ow_carry(w_carry_26_26));
wire w_sum_26_24, w_carry_26_24;
math_adder_full FA_26_24(.i_a(w_carry_25_20), .i_b(w_carry_25_18), .i_c(w_carry_25_16), .ow_sum(w_sum_26_24), .ow_carry(w_carry_26_24));
wire w_sum_26_22, w_carry_26_22;
math_adder_full FA_26_22(.i_a(w_carry_25_14), .i_b(w_carry_25_12), .i_c(w_carry_25_10), .ow_sum(w_sum_26_22), .ow_carry(w_carry_26_22));
wire w_sum_26_20, w_carry_26_20;
math_adder_full FA_26_20(.i_a(w_carry_25_08), .i_b(w_carry_25_06), .i_c(w_carry_25_04), .ow_sum(w_sum_26_20), .ow_carry(w_carry_26_20));
wire w_sum_26_18, w_carry_26_18;
math_adder_full FA_26_18(.i_a(w_carry_25_02), .i_b(w_sum_26_52), .i_c(w_sum_26_50), .ow_sum(w_sum_26_18), .ow_carry(w_carry_26_18));
wire w_sum_26_16, w_carry_26_16;
math_adder_full FA_26_16(.i_a(w_sum_26_48), .i_b(w_sum_26_46), .i_c(w_sum_26_44), .ow_sum(w_sum_26_16), .ow_carry(w_carry_26_16));
wire w_sum_26_14, w_carry_26_14;
math_adder_full FA_26_14(.i_a(w_sum_26_42), .i_b(w_sum_26_40), .i_c(w_sum_26_38), .ow_sum(w_sum_26_14), .ow_carry(w_carry_26_14));
wire w_sum_26_12, w_carry_26_12;
math_adder_full FA_26_12(.i_a(w_sum_26_36), .i_b(w_sum_26_34), .i_c(w_sum_26_32), .ow_sum(w_sum_26_12), .ow_carry(w_carry_26_12));
wire w_sum_26_10, w_carry_26_10;
math_adder_full FA_26_10(.i_a(w_sum_26_30), .i_b(w_sum_26_28), .i_c(w_sum_26_26), .ow_sum(w_sum_26_10), .ow_carry(w_carry_26_10));
wire w_sum_26_08, w_carry_26_08;
math_adder_full FA_26_08(.i_a(w_sum_26_24), .i_b(w_sum_26_22), .i_c(w_sum_26_20), .ow_sum(w_sum_26_08), .ow_carry(w_carry_26_08));
wire w_sum_26_06, w_carry_26_06;
math_adder_full FA_26_06(.i_a(w_sum_26_18), .i_b(w_sum_26_16), .i_c(w_sum_26_14), .ow_sum(w_sum_26_06), .ow_carry(w_carry_26_06));
wire w_sum_26_04, w_carry_26_04;
math_adder_full FA_26_04(.i_a(w_sum_26_12), .i_b(w_sum_26_10), .i_c(w_sum_26_08), .ow_sum(w_sum_26_04), .ow_carry(w_carry_26_04));
wire w_sum_26_02, w_carry_26_02;
math_adder_half HA_26_02(.i_a(w_sum_26_06), .i_b(w_sum_26_04), .ow_sum(w_sum_26_02), .ow_carry(w_carry_26_02));
wire w_sum_27_54, w_carry_27_54;
math_adder_full FA_27_54(.i_a(w_pp_00_27), .i_b(w_pp_01_26), .i_c(w_pp_02_25), .ow_sum(w_sum_27_54), .ow_carry(w_carry_27_54));
wire w_sum_27_52, w_carry_27_52;
math_adder_full FA_27_52(.i_a(w_pp_03_24), .i_b(w_pp_04_23), .i_c(w_pp_05_22), .ow_sum(w_sum_27_52), .ow_carry(w_carry_27_52));
wire w_sum_27_50, w_carry_27_50;
math_adder_full FA_27_50(.i_a(w_pp_06_21), .i_b(w_pp_07_20), .i_c(w_pp_08_19), .ow_sum(w_sum_27_50), .ow_carry(w_carry_27_50));
wire w_sum_27_48, w_carry_27_48;
math_adder_full FA_27_48(.i_a(w_pp_09_18), .i_b(w_pp_10_17), .i_c(w_pp_11_16), .ow_sum(w_sum_27_48), .ow_carry(w_carry_27_48));
wire w_sum_27_46, w_carry_27_46;
math_adder_full FA_27_46(.i_a(w_pp_12_15), .i_b(w_pp_13_14), .i_c(w_pp_14_13), .ow_sum(w_sum_27_46), .ow_carry(w_carry_27_46));
wire w_sum_27_44, w_carry_27_44;
math_adder_full FA_27_44(.i_a(w_pp_15_12), .i_b(w_pp_16_11), .i_c(w_pp_17_10), .ow_sum(w_sum_27_44), .ow_carry(w_carry_27_44));
wire w_sum_27_42, w_carry_27_42;
math_adder_full FA_27_42(.i_a(w_pp_18_09), .i_b(w_pp_19_08), .i_c(w_pp_20_07), .ow_sum(w_sum_27_42), .ow_carry(w_carry_27_42));
wire w_sum_27_40, w_carry_27_40;
math_adder_full FA_27_40(.i_a(w_pp_21_06), .i_b(w_pp_22_05), .i_c(w_pp_23_04), .ow_sum(w_sum_27_40), .ow_carry(w_carry_27_40));
wire w_sum_27_38, w_carry_27_38;
math_adder_full FA_27_38(.i_a(w_pp_24_03), .i_b(w_pp_25_02), .i_c(w_pp_26_01), .ow_sum(w_sum_27_38), .ow_carry(w_carry_27_38));
wire w_sum_27_36, w_carry_27_36;
math_adder_full FA_27_36(.i_a(w_pp_27_00), .i_b(w_carry_26_52), .i_c(w_carry_26_50), .ow_sum(w_sum_27_36), .ow_carry(w_carry_27_36));
wire w_sum_27_34, w_carry_27_34;
math_adder_full FA_27_34(.i_a(w_carry_26_48), .i_b(w_carry_26_46), .i_c(w_carry_26_44), .ow_sum(w_sum_27_34), .ow_carry(w_carry_27_34));
wire w_sum_27_32, w_carry_27_32;
math_adder_full FA_27_32(.i_a(w_carry_26_42), .i_b(w_carry_26_40), .i_c(w_carry_26_38), .ow_sum(w_sum_27_32), .ow_carry(w_carry_27_32));
wire w_sum_27_30, w_carry_27_30;
math_adder_full FA_27_30(.i_a(w_carry_26_36), .i_b(w_carry_26_34), .i_c(w_carry_26_32), .ow_sum(w_sum_27_30), .ow_carry(w_carry_27_30));
wire w_sum_27_28, w_carry_27_28;
math_adder_full FA_27_28(.i_a(w_carry_26_30), .i_b(w_carry_26_28), .i_c(w_carry_26_26), .ow_sum(w_sum_27_28), .ow_carry(w_carry_27_28));
wire w_sum_27_26, w_carry_27_26;
math_adder_full FA_27_26(.i_a(w_carry_26_24), .i_b(w_carry_26_22), .i_c(w_carry_26_20), .ow_sum(w_sum_27_26), .ow_carry(w_carry_27_26));
wire w_sum_27_24, w_carry_27_24;
math_adder_full FA_27_24(.i_a(w_carry_26_18), .i_b(w_carry_26_16), .i_c(w_carry_26_14), .ow_sum(w_sum_27_24), .ow_carry(w_carry_27_24));
wire w_sum_27_22, w_carry_27_22;
math_adder_full FA_27_22(.i_a(w_carry_26_12), .i_b(w_carry_26_10), .i_c(w_carry_26_08), .ow_sum(w_sum_27_22), .ow_carry(w_carry_27_22));
wire w_sum_27_20, w_carry_27_20;
math_adder_full FA_27_20(.i_a(w_carry_26_06), .i_b(w_carry_26_04), .i_c(w_carry_26_02), .ow_sum(w_sum_27_20), .ow_carry(w_carry_27_20));
wire w_sum_27_18, w_carry_27_18;
math_adder_full FA_27_18(.i_a(w_sum_27_54), .i_b(w_sum_27_52), .i_c(w_sum_27_50), .ow_sum(w_sum_27_18), .ow_carry(w_carry_27_18));
wire w_sum_27_16, w_carry_27_16;
math_adder_full FA_27_16(.i_a(w_sum_27_48), .i_b(w_sum_27_46), .i_c(w_sum_27_44), .ow_sum(w_sum_27_16), .ow_carry(w_carry_27_16));
wire w_sum_27_14, w_carry_27_14;
math_adder_full FA_27_14(.i_a(w_sum_27_42), .i_b(w_sum_27_40), .i_c(w_sum_27_38), .ow_sum(w_sum_27_14), .ow_carry(w_carry_27_14));
wire w_sum_27_12, w_carry_27_12;
math_adder_full FA_27_12(.i_a(w_sum_27_36), .i_b(w_sum_27_34), .i_c(w_sum_27_32), .ow_sum(w_sum_27_12), .ow_carry(w_carry_27_12));
wire w_sum_27_10, w_carry_27_10;
math_adder_full FA_27_10(.i_a(w_sum_27_30), .i_b(w_sum_27_28), .i_c(w_sum_27_26), .ow_sum(w_sum_27_10), .ow_carry(w_carry_27_10));
wire w_sum_27_08, w_carry_27_08;
math_adder_full FA_27_08(.i_a(w_sum_27_24), .i_b(w_sum_27_22), .i_c(w_sum_27_20), .ow_sum(w_sum_27_08), .ow_carry(w_carry_27_08));
wire w_sum_27_06, w_carry_27_06;
math_adder_full FA_27_06(.i_a(w_sum_27_18), .i_b(w_sum_27_16), .i_c(w_sum_27_14), .ow_sum(w_sum_27_06), .ow_carry(w_carry_27_06));
wire w_sum_27_04, w_carry_27_04;
math_adder_full FA_27_04(.i_a(w_sum_27_12), .i_b(w_sum_27_10), .i_c(w_sum_27_08), .ow_sum(w_sum_27_04), .ow_carry(w_carry_27_04));
wire w_sum_27_02, w_carry_27_02;
math_adder_half HA_27_02(.i_a(w_sum_27_06), .i_b(w_sum_27_04), .ow_sum(w_sum_27_02), .ow_carry(w_carry_27_02));
wire w_sum_28_56, w_carry_28_56;
math_adder_full FA_28_56(.i_a(w_pp_00_28), .i_b(w_pp_01_27), .i_c(w_pp_02_26), .ow_sum(w_sum_28_56), .ow_carry(w_carry_28_56));
wire w_sum_28_54, w_carry_28_54;
math_adder_full FA_28_54(.i_a(w_pp_03_25), .i_b(w_pp_04_24), .i_c(w_pp_05_23), .ow_sum(w_sum_28_54), .ow_carry(w_carry_28_54));
wire w_sum_28_52, w_carry_28_52;
math_adder_full FA_28_52(.i_a(w_pp_06_22), .i_b(w_pp_07_21), .i_c(w_pp_08_20), .ow_sum(w_sum_28_52), .ow_carry(w_carry_28_52));
wire w_sum_28_50, w_carry_28_50;
math_adder_full FA_28_50(.i_a(w_pp_09_19), .i_b(w_pp_10_18), .i_c(w_pp_11_17), .ow_sum(w_sum_28_50), .ow_carry(w_carry_28_50));
wire w_sum_28_48, w_carry_28_48;
math_adder_full FA_28_48(.i_a(w_pp_12_16), .i_b(w_pp_13_15), .i_c(w_pp_14_14), .ow_sum(w_sum_28_48), .ow_carry(w_carry_28_48));
wire w_sum_28_46, w_carry_28_46;
math_adder_full FA_28_46(.i_a(w_pp_15_13), .i_b(w_pp_16_12), .i_c(w_pp_17_11), .ow_sum(w_sum_28_46), .ow_carry(w_carry_28_46));
wire w_sum_28_44, w_carry_28_44;
math_adder_full FA_28_44(.i_a(w_pp_18_10), .i_b(w_pp_19_09), .i_c(w_pp_20_08), .ow_sum(w_sum_28_44), .ow_carry(w_carry_28_44));
wire w_sum_28_42, w_carry_28_42;
math_adder_full FA_28_42(.i_a(w_pp_21_07), .i_b(w_pp_22_06), .i_c(w_pp_23_05), .ow_sum(w_sum_28_42), .ow_carry(w_carry_28_42));
wire w_sum_28_40, w_carry_28_40;
math_adder_full FA_28_40(.i_a(w_pp_24_04), .i_b(w_pp_25_03), .i_c(w_pp_26_02), .ow_sum(w_sum_28_40), .ow_carry(w_carry_28_40));
wire w_sum_28_38, w_carry_28_38;
math_adder_full FA_28_38(.i_a(w_pp_27_01), .i_b(w_pp_28_00), .i_c(w_carry_27_54), .ow_sum(w_sum_28_38), .ow_carry(w_carry_28_38));
wire w_sum_28_36, w_carry_28_36;
math_adder_full FA_28_36(.i_a(w_carry_27_52), .i_b(w_carry_27_50), .i_c(w_carry_27_48), .ow_sum(w_sum_28_36), .ow_carry(w_carry_28_36));
wire w_sum_28_34, w_carry_28_34;
math_adder_full FA_28_34(.i_a(w_carry_27_46), .i_b(w_carry_27_44), .i_c(w_carry_27_42), .ow_sum(w_sum_28_34), .ow_carry(w_carry_28_34));
wire w_sum_28_32, w_carry_28_32;
math_adder_full FA_28_32(.i_a(w_carry_27_40), .i_b(w_carry_27_38), .i_c(w_carry_27_36), .ow_sum(w_sum_28_32), .ow_carry(w_carry_28_32));
wire w_sum_28_30, w_carry_28_30;
math_adder_full FA_28_30(.i_a(w_carry_27_34), .i_b(w_carry_27_32), .i_c(w_carry_27_30), .ow_sum(w_sum_28_30), .ow_carry(w_carry_28_30));
wire w_sum_28_28, w_carry_28_28;
math_adder_full FA_28_28(.i_a(w_carry_27_28), .i_b(w_carry_27_26), .i_c(w_carry_27_24), .ow_sum(w_sum_28_28), .ow_carry(w_carry_28_28));
wire w_sum_28_26, w_carry_28_26;
math_adder_full FA_28_26(.i_a(w_carry_27_22), .i_b(w_carry_27_20), .i_c(w_carry_27_18), .ow_sum(w_sum_28_26), .ow_carry(w_carry_28_26));
wire w_sum_28_24, w_carry_28_24;
math_adder_full FA_28_24(.i_a(w_carry_27_16), .i_b(w_carry_27_14), .i_c(w_carry_27_12), .ow_sum(w_sum_28_24), .ow_carry(w_carry_28_24));
wire w_sum_28_22, w_carry_28_22;
math_adder_full FA_28_22(.i_a(w_carry_27_10), .i_b(w_carry_27_08), .i_c(w_carry_27_06), .ow_sum(w_sum_28_22), .ow_carry(w_carry_28_22));
wire w_sum_28_20, w_carry_28_20;
math_adder_full FA_28_20(.i_a(w_carry_27_04), .i_b(w_carry_27_02), .i_c(w_sum_28_56), .ow_sum(w_sum_28_20), .ow_carry(w_carry_28_20));
wire w_sum_28_18, w_carry_28_18;
math_adder_full FA_28_18(.i_a(w_sum_28_54), .i_b(w_sum_28_52), .i_c(w_sum_28_50), .ow_sum(w_sum_28_18), .ow_carry(w_carry_28_18));
wire w_sum_28_16, w_carry_28_16;
math_adder_full FA_28_16(.i_a(w_sum_28_48), .i_b(w_sum_28_46), .i_c(w_sum_28_44), .ow_sum(w_sum_28_16), .ow_carry(w_carry_28_16));
wire w_sum_28_14, w_carry_28_14;
math_adder_full FA_28_14(.i_a(w_sum_28_42), .i_b(w_sum_28_40), .i_c(w_sum_28_38), .ow_sum(w_sum_28_14), .ow_carry(w_carry_28_14));
wire w_sum_28_12, w_carry_28_12;
math_adder_full FA_28_12(.i_a(w_sum_28_36), .i_b(w_sum_28_34), .i_c(w_sum_28_32), .ow_sum(w_sum_28_12), .ow_carry(w_carry_28_12));
wire w_sum_28_10, w_carry_28_10;
math_adder_full FA_28_10(.i_a(w_sum_28_30), .i_b(w_sum_28_28), .i_c(w_sum_28_26), .ow_sum(w_sum_28_10), .ow_carry(w_carry_28_10));
wire w_sum_28_08, w_carry_28_08;
math_adder_full FA_28_08(.i_a(w_sum_28_24), .i_b(w_sum_28_22), .i_c(w_sum_28_20), .ow_sum(w_sum_28_08), .ow_carry(w_carry_28_08));
wire w_sum_28_06, w_carry_28_06;
math_adder_full FA_28_06(.i_a(w_sum_28_18), .i_b(w_sum_28_16), .i_c(w_sum_28_14), .ow_sum(w_sum_28_06), .ow_carry(w_carry_28_06));
wire w_sum_28_04, w_carry_28_04;
math_adder_full FA_28_04(.i_a(w_sum_28_12), .i_b(w_sum_28_10), .i_c(w_sum_28_08), .ow_sum(w_sum_28_04), .ow_carry(w_carry_28_04));
wire w_sum_28_02, w_carry_28_02;
math_adder_half HA_28_02(.i_a(w_sum_28_06), .i_b(w_sum_28_04), .ow_sum(w_sum_28_02), .ow_carry(w_carry_28_02));
wire w_sum_29_58, w_carry_29_58;
math_adder_full FA_29_58(.i_a(w_pp_00_29), .i_b(w_pp_01_28), .i_c(w_pp_02_27), .ow_sum(w_sum_29_58), .ow_carry(w_carry_29_58));
wire w_sum_29_56, w_carry_29_56;
math_adder_full FA_29_56(.i_a(w_pp_03_26), .i_b(w_pp_04_25), .i_c(w_pp_05_24), .ow_sum(w_sum_29_56), .ow_carry(w_carry_29_56));
wire w_sum_29_54, w_carry_29_54;
math_adder_full FA_29_54(.i_a(w_pp_06_23), .i_b(w_pp_07_22), .i_c(w_pp_08_21), .ow_sum(w_sum_29_54), .ow_carry(w_carry_29_54));
wire w_sum_29_52, w_carry_29_52;
math_adder_full FA_29_52(.i_a(w_pp_09_20), .i_b(w_pp_10_19), .i_c(w_pp_11_18), .ow_sum(w_sum_29_52), .ow_carry(w_carry_29_52));
wire w_sum_29_50, w_carry_29_50;
math_adder_full FA_29_50(.i_a(w_pp_12_17), .i_b(w_pp_13_16), .i_c(w_pp_14_15), .ow_sum(w_sum_29_50), .ow_carry(w_carry_29_50));
wire w_sum_29_48, w_carry_29_48;
math_adder_full FA_29_48(.i_a(w_pp_15_14), .i_b(w_pp_16_13), .i_c(w_pp_17_12), .ow_sum(w_sum_29_48), .ow_carry(w_carry_29_48));
wire w_sum_29_46, w_carry_29_46;
math_adder_full FA_29_46(.i_a(w_pp_18_11), .i_b(w_pp_19_10), .i_c(w_pp_20_09), .ow_sum(w_sum_29_46), .ow_carry(w_carry_29_46));
wire w_sum_29_44, w_carry_29_44;
math_adder_full FA_29_44(.i_a(w_pp_21_08), .i_b(w_pp_22_07), .i_c(w_pp_23_06), .ow_sum(w_sum_29_44), .ow_carry(w_carry_29_44));
wire w_sum_29_42, w_carry_29_42;
math_adder_full FA_29_42(.i_a(w_pp_24_05), .i_b(w_pp_25_04), .i_c(w_pp_26_03), .ow_sum(w_sum_29_42), .ow_carry(w_carry_29_42));
wire w_sum_29_40, w_carry_29_40;
math_adder_full FA_29_40(.i_a(w_pp_27_02), .i_b(w_pp_28_01), .i_c(w_pp_29_00), .ow_sum(w_sum_29_40), .ow_carry(w_carry_29_40));
wire w_sum_29_38, w_carry_29_38;
math_adder_full FA_29_38(.i_a(w_carry_28_56), .i_b(w_carry_28_54), .i_c(w_carry_28_52), .ow_sum(w_sum_29_38), .ow_carry(w_carry_29_38));
wire w_sum_29_36, w_carry_29_36;
math_adder_full FA_29_36(.i_a(w_carry_28_50), .i_b(w_carry_28_48), .i_c(w_carry_28_46), .ow_sum(w_sum_29_36), .ow_carry(w_carry_29_36));
wire w_sum_29_34, w_carry_29_34;
math_adder_full FA_29_34(.i_a(w_carry_28_44), .i_b(w_carry_28_42), .i_c(w_carry_28_40), .ow_sum(w_sum_29_34), .ow_carry(w_carry_29_34));
wire w_sum_29_32, w_carry_29_32;
math_adder_full FA_29_32(.i_a(w_carry_28_38), .i_b(w_carry_28_36), .i_c(w_carry_28_34), .ow_sum(w_sum_29_32), .ow_carry(w_carry_29_32));
wire w_sum_29_30, w_carry_29_30;
math_adder_full FA_29_30(.i_a(w_carry_28_32), .i_b(w_carry_28_30), .i_c(w_carry_28_28), .ow_sum(w_sum_29_30), .ow_carry(w_carry_29_30));
wire w_sum_29_28, w_carry_29_28;
math_adder_full FA_29_28(.i_a(w_carry_28_26), .i_b(w_carry_28_24), .i_c(w_carry_28_22), .ow_sum(w_sum_29_28), .ow_carry(w_carry_29_28));
wire w_sum_29_26, w_carry_29_26;
math_adder_full FA_29_26(.i_a(w_carry_28_20), .i_b(w_carry_28_18), .i_c(w_carry_28_16), .ow_sum(w_sum_29_26), .ow_carry(w_carry_29_26));
wire w_sum_29_24, w_carry_29_24;
math_adder_full FA_29_24(.i_a(w_carry_28_14), .i_b(w_carry_28_12), .i_c(w_carry_28_10), .ow_sum(w_sum_29_24), .ow_carry(w_carry_29_24));
wire w_sum_29_22, w_carry_29_22;
math_adder_full FA_29_22(.i_a(w_carry_28_08), .i_b(w_carry_28_06), .i_c(w_carry_28_04), .ow_sum(w_sum_29_22), .ow_carry(w_carry_29_22));
wire w_sum_29_20, w_carry_29_20;
math_adder_full FA_29_20(.i_a(w_carry_28_02), .i_b(w_sum_29_58), .i_c(w_sum_29_56), .ow_sum(w_sum_29_20), .ow_carry(w_carry_29_20));
wire w_sum_29_18, w_carry_29_18;
math_adder_full FA_29_18(.i_a(w_sum_29_54), .i_b(w_sum_29_52), .i_c(w_sum_29_50), .ow_sum(w_sum_29_18), .ow_carry(w_carry_29_18));
wire w_sum_29_16, w_carry_29_16;
math_adder_full FA_29_16(.i_a(w_sum_29_48), .i_b(w_sum_29_46), .i_c(w_sum_29_44), .ow_sum(w_sum_29_16), .ow_carry(w_carry_29_16));
wire w_sum_29_14, w_carry_29_14;
math_adder_full FA_29_14(.i_a(w_sum_29_42), .i_b(w_sum_29_40), .i_c(w_sum_29_38), .ow_sum(w_sum_29_14), .ow_carry(w_carry_29_14));
wire w_sum_29_12, w_carry_29_12;
math_adder_full FA_29_12(.i_a(w_sum_29_36), .i_b(w_sum_29_34), .i_c(w_sum_29_32), .ow_sum(w_sum_29_12), .ow_carry(w_carry_29_12));
wire w_sum_29_10, w_carry_29_10;
math_adder_full FA_29_10(.i_a(w_sum_29_30), .i_b(w_sum_29_28), .i_c(w_sum_29_26), .ow_sum(w_sum_29_10), .ow_carry(w_carry_29_10));
wire w_sum_29_08, w_carry_29_08;
math_adder_full FA_29_08(.i_a(w_sum_29_24), .i_b(w_sum_29_22), .i_c(w_sum_29_20), .ow_sum(w_sum_29_08), .ow_carry(w_carry_29_08));
wire w_sum_29_06, w_carry_29_06;
math_adder_full FA_29_06(.i_a(w_sum_29_18), .i_b(w_sum_29_16), .i_c(w_sum_29_14), .ow_sum(w_sum_29_06), .ow_carry(w_carry_29_06));
wire w_sum_29_04, w_carry_29_04;
math_adder_full FA_29_04(.i_a(w_sum_29_12), .i_b(w_sum_29_10), .i_c(w_sum_29_08), .ow_sum(w_sum_29_04), .ow_carry(w_carry_29_04));
wire w_sum_29_02, w_carry_29_02;
math_adder_half HA_29_02(.i_a(w_sum_29_06), .i_b(w_sum_29_04), .ow_sum(w_sum_29_02), .ow_carry(w_carry_29_02));
wire w_sum_30_60, w_carry_30_60;
math_adder_full FA_30_60(.i_a(w_pp_00_30), .i_b(w_pp_01_29), .i_c(w_pp_02_28), .ow_sum(w_sum_30_60), .ow_carry(w_carry_30_60));
wire w_sum_30_58, w_carry_30_58;
math_adder_full FA_30_58(.i_a(w_pp_03_27), .i_b(w_pp_04_26), .i_c(w_pp_05_25), .ow_sum(w_sum_30_58), .ow_carry(w_carry_30_58));
wire w_sum_30_56, w_carry_30_56;
math_adder_full FA_30_56(.i_a(w_pp_06_24), .i_b(w_pp_07_23), .i_c(w_pp_08_22), .ow_sum(w_sum_30_56), .ow_carry(w_carry_30_56));
wire w_sum_30_54, w_carry_30_54;
math_adder_full FA_30_54(.i_a(w_pp_09_21), .i_b(w_pp_10_20), .i_c(w_pp_11_19), .ow_sum(w_sum_30_54), .ow_carry(w_carry_30_54));
wire w_sum_30_52, w_carry_30_52;
math_adder_full FA_30_52(.i_a(w_pp_12_18), .i_b(w_pp_13_17), .i_c(w_pp_14_16), .ow_sum(w_sum_30_52), .ow_carry(w_carry_30_52));
wire w_sum_30_50, w_carry_30_50;
math_adder_full FA_30_50(.i_a(w_pp_15_15), .i_b(w_pp_16_14), .i_c(w_pp_17_13), .ow_sum(w_sum_30_50), .ow_carry(w_carry_30_50));
wire w_sum_30_48, w_carry_30_48;
math_adder_full FA_30_48(.i_a(w_pp_18_12), .i_b(w_pp_19_11), .i_c(w_pp_20_10), .ow_sum(w_sum_30_48), .ow_carry(w_carry_30_48));
wire w_sum_30_46, w_carry_30_46;
math_adder_full FA_30_46(.i_a(w_pp_21_09), .i_b(w_pp_22_08), .i_c(w_pp_23_07), .ow_sum(w_sum_30_46), .ow_carry(w_carry_30_46));
wire w_sum_30_44, w_carry_30_44;
math_adder_full FA_30_44(.i_a(w_pp_24_06), .i_b(w_pp_25_05), .i_c(w_pp_26_04), .ow_sum(w_sum_30_44), .ow_carry(w_carry_30_44));
wire w_sum_30_42, w_carry_30_42;
math_adder_full FA_30_42(.i_a(w_pp_27_03), .i_b(w_pp_28_02), .i_c(w_pp_29_01), .ow_sum(w_sum_30_42), .ow_carry(w_carry_30_42));
wire w_sum_30_40, w_carry_30_40;
math_adder_full FA_30_40(.i_a(w_pp_30_00), .i_b(w_carry_29_58), .i_c(w_carry_29_56), .ow_sum(w_sum_30_40), .ow_carry(w_carry_30_40));
wire w_sum_30_38, w_carry_30_38;
math_adder_full FA_30_38(.i_a(w_carry_29_54), .i_b(w_carry_29_52), .i_c(w_carry_29_50), .ow_sum(w_sum_30_38), .ow_carry(w_carry_30_38));
wire w_sum_30_36, w_carry_30_36;
math_adder_full FA_30_36(.i_a(w_carry_29_48), .i_b(w_carry_29_46), .i_c(w_carry_29_44), .ow_sum(w_sum_30_36), .ow_carry(w_carry_30_36));
wire w_sum_30_34, w_carry_30_34;
math_adder_full FA_30_34(.i_a(w_carry_29_42), .i_b(w_carry_29_40), .i_c(w_carry_29_38), .ow_sum(w_sum_30_34), .ow_carry(w_carry_30_34));
wire w_sum_30_32, w_carry_30_32;
math_adder_full FA_30_32(.i_a(w_carry_29_36), .i_b(w_carry_29_34), .i_c(w_carry_29_32), .ow_sum(w_sum_30_32), .ow_carry(w_carry_30_32));
wire w_sum_30_30, w_carry_30_30;
math_adder_full FA_30_30(.i_a(w_carry_29_30), .i_b(w_carry_29_28), .i_c(w_carry_29_26), .ow_sum(w_sum_30_30), .ow_carry(w_carry_30_30));
wire w_sum_30_28, w_carry_30_28;
math_adder_full FA_30_28(.i_a(w_carry_29_24), .i_b(w_carry_29_22), .i_c(w_carry_29_20), .ow_sum(w_sum_30_28), .ow_carry(w_carry_30_28));
wire w_sum_30_26, w_carry_30_26;
math_adder_full FA_30_26(.i_a(w_carry_29_18), .i_b(w_carry_29_16), .i_c(w_carry_29_14), .ow_sum(w_sum_30_26), .ow_carry(w_carry_30_26));
wire w_sum_30_24, w_carry_30_24;
math_adder_full FA_30_24(.i_a(w_carry_29_12), .i_b(w_carry_29_10), .i_c(w_carry_29_08), .ow_sum(w_sum_30_24), .ow_carry(w_carry_30_24));
wire w_sum_30_22, w_carry_30_22;
math_adder_full FA_30_22(.i_a(w_carry_29_06), .i_b(w_carry_29_04), .i_c(w_carry_29_02), .ow_sum(w_sum_30_22), .ow_carry(w_carry_30_22));
wire w_sum_30_20, w_carry_30_20;
math_adder_full FA_30_20(.i_a(w_sum_30_60), .i_b(w_sum_30_58), .i_c(w_sum_30_56), .ow_sum(w_sum_30_20), .ow_carry(w_carry_30_20));
wire w_sum_30_18, w_carry_30_18;
math_adder_full FA_30_18(.i_a(w_sum_30_54), .i_b(w_sum_30_52), .i_c(w_sum_30_50), .ow_sum(w_sum_30_18), .ow_carry(w_carry_30_18));
wire w_sum_30_16, w_carry_30_16;
math_adder_full FA_30_16(.i_a(w_sum_30_48), .i_b(w_sum_30_46), .i_c(w_sum_30_44), .ow_sum(w_sum_30_16), .ow_carry(w_carry_30_16));
wire w_sum_30_14, w_carry_30_14;
math_adder_full FA_30_14(.i_a(w_sum_30_42), .i_b(w_sum_30_40), .i_c(w_sum_30_38), .ow_sum(w_sum_30_14), .ow_carry(w_carry_30_14));
wire w_sum_30_12, w_carry_30_12;
math_adder_full FA_30_12(.i_a(w_sum_30_36), .i_b(w_sum_30_34), .i_c(w_sum_30_32), .ow_sum(w_sum_30_12), .ow_carry(w_carry_30_12));
wire w_sum_30_10, w_carry_30_10;
math_adder_full FA_30_10(.i_a(w_sum_30_30), .i_b(w_sum_30_28), .i_c(w_sum_30_26), .ow_sum(w_sum_30_10), .ow_carry(w_carry_30_10));
wire w_sum_30_08, w_carry_30_08;
math_adder_full FA_30_08(.i_a(w_sum_30_24), .i_b(w_sum_30_22), .i_c(w_sum_30_20), .ow_sum(w_sum_30_08), .ow_carry(w_carry_30_08));
wire w_sum_30_06, w_carry_30_06;
math_adder_full FA_30_06(.i_a(w_sum_30_18), .i_b(w_sum_30_16), .i_c(w_sum_30_14), .ow_sum(w_sum_30_06), .ow_carry(w_carry_30_06));
wire w_sum_30_04, w_carry_30_04;
math_adder_full FA_30_04(.i_a(w_sum_30_12), .i_b(w_sum_30_10), .i_c(w_sum_30_08), .ow_sum(w_sum_30_04), .ow_carry(w_carry_30_04));
wire w_sum_30_02, w_carry_30_02;
math_adder_half HA_30_02(.i_a(w_sum_30_06), .i_b(w_sum_30_04), .ow_sum(w_sum_30_02), .ow_carry(w_carry_30_02));
wire w_sum_31_62, w_carry_31_62;
math_adder_full FA_31_62(.i_a(w_pp_00_31), .i_b(w_pp_01_30), .i_c(w_pp_02_29), .ow_sum(w_sum_31_62), .ow_carry(w_carry_31_62));
wire w_sum_31_60, w_carry_31_60;
math_adder_full FA_31_60(.i_a(w_pp_03_28), .i_b(w_pp_04_27), .i_c(w_pp_05_26), .ow_sum(w_sum_31_60), .ow_carry(w_carry_31_60));
wire w_sum_31_58, w_carry_31_58;
math_adder_full FA_31_58(.i_a(w_pp_06_25), .i_b(w_pp_07_24), .i_c(w_pp_08_23), .ow_sum(w_sum_31_58), .ow_carry(w_carry_31_58));
wire w_sum_31_56, w_carry_31_56;
math_adder_full FA_31_56(.i_a(w_pp_09_22), .i_b(w_pp_10_21), .i_c(w_pp_11_20), .ow_sum(w_sum_31_56), .ow_carry(w_carry_31_56));
wire w_sum_31_54, w_carry_31_54;
math_adder_full FA_31_54(.i_a(w_pp_12_19), .i_b(w_pp_13_18), .i_c(w_pp_14_17), .ow_sum(w_sum_31_54), .ow_carry(w_carry_31_54));
wire w_sum_31_52, w_carry_31_52;
math_adder_full FA_31_52(.i_a(w_pp_15_16), .i_b(w_pp_16_15), .i_c(w_pp_17_14), .ow_sum(w_sum_31_52), .ow_carry(w_carry_31_52));
wire w_sum_31_50, w_carry_31_50;
math_adder_full FA_31_50(.i_a(w_pp_18_13), .i_b(w_pp_19_12), .i_c(w_pp_20_11), .ow_sum(w_sum_31_50), .ow_carry(w_carry_31_50));
wire w_sum_31_48, w_carry_31_48;
math_adder_full FA_31_48(.i_a(w_pp_21_10), .i_b(w_pp_22_09), .i_c(w_pp_23_08), .ow_sum(w_sum_31_48), .ow_carry(w_carry_31_48));
wire w_sum_31_46, w_carry_31_46;
math_adder_full FA_31_46(.i_a(w_pp_24_07), .i_b(w_pp_25_06), .i_c(w_pp_26_05), .ow_sum(w_sum_31_46), .ow_carry(w_carry_31_46));
wire w_sum_31_44, w_carry_31_44;
math_adder_full FA_31_44(.i_a(w_pp_27_04), .i_b(w_pp_28_03), .i_c(w_pp_29_02), .ow_sum(w_sum_31_44), .ow_carry(w_carry_31_44));
wire w_sum_31_42, w_carry_31_42;
math_adder_full FA_31_42(.i_a(w_pp_30_01), .i_b(w_pp_31_00), .i_c(w_carry_30_60), .ow_sum(w_sum_31_42), .ow_carry(w_carry_31_42));
wire w_sum_31_40, w_carry_31_40;
math_adder_full FA_31_40(.i_a(w_carry_30_58), .i_b(w_carry_30_56), .i_c(w_carry_30_54), .ow_sum(w_sum_31_40), .ow_carry(w_carry_31_40));
wire w_sum_31_38, w_carry_31_38;
math_adder_full FA_31_38(.i_a(w_carry_30_52), .i_b(w_carry_30_50), .i_c(w_carry_30_48), .ow_sum(w_sum_31_38), .ow_carry(w_carry_31_38));
wire w_sum_31_36, w_carry_31_36;
math_adder_full FA_31_36(.i_a(w_carry_30_46), .i_b(w_carry_30_44), .i_c(w_carry_30_42), .ow_sum(w_sum_31_36), .ow_carry(w_carry_31_36));
wire w_sum_31_34, w_carry_31_34;
math_adder_full FA_31_34(.i_a(w_carry_30_40), .i_b(w_carry_30_38), .i_c(w_carry_30_36), .ow_sum(w_sum_31_34), .ow_carry(w_carry_31_34));
wire w_sum_31_32, w_carry_31_32;
math_adder_full FA_31_32(.i_a(w_carry_30_34), .i_b(w_carry_30_32), .i_c(w_carry_30_30), .ow_sum(w_sum_31_32), .ow_carry(w_carry_31_32));
wire w_sum_31_30, w_carry_31_30;
math_adder_full FA_31_30(.i_a(w_carry_30_28), .i_b(w_carry_30_26), .i_c(w_carry_30_24), .ow_sum(w_sum_31_30), .ow_carry(w_carry_31_30));
wire w_sum_31_28, w_carry_31_28;
math_adder_full FA_31_28(.i_a(w_carry_30_22), .i_b(w_carry_30_20), .i_c(w_carry_30_18), .ow_sum(w_sum_31_28), .ow_carry(w_carry_31_28));
wire w_sum_31_26, w_carry_31_26;
math_adder_full FA_31_26(.i_a(w_carry_30_16), .i_b(w_carry_30_14), .i_c(w_carry_30_12), .ow_sum(w_sum_31_26), .ow_carry(w_carry_31_26));
wire w_sum_31_24, w_carry_31_24;
math_adder_full FA_31_24(.i_a(w_carry_30_10), .i_b(w_carry_30_08), .i_c(w_carry_30_06), .ow_sum(w_sum_31_24), .ow_carry(w_carry_31_24));
wire w_sum_31_22, w_carry_31_22;
math_adder_full FA_31_22(.i_a(w_carry_30_04), .i_b(w_carry_30_02), .i_c(w_sum_31_62), .ow_sum(w_sum_31_22), .ow_carry(w_carry_31_22));
wire w_sum_31_20, w_carry_31_20;
math_adder_full FA_31_20(.i_a(w_sum_31_60), .i_b(w_sum_31_58), .i_c(w_sum_31_56), .ow_sum(w_sum_31_20), .ow_carry(w_carry_31_20));
wire w_sum_31_18, w_carry_31_18;
math_adder_full FA_31_18(.i_a(w_sum_31_54), .i_b(w_sum_31_52), .i_c(w_sum_31_50), .ow_sum(w_sum_31_18), .ow_carry(w_carry_31_18));
wire w_sum_31_16, w_carry_31_16;
math_adder_full FA_31_16(.i_a(w_sum_31_48), .i_b(w_sum_31_46), .i_c(w_sum_31_44), .ow_sum(w_sum_31_16), .ow_carry(w_carry_31_16));
wire w_sum_31_14, w_carry_31_14;
math_adder_full FA_31_14(.i_a(w_sum_31_42), .i_b(w_sum_31_40), .i_c(w_sum_31_38), .ow_sum(w_sum_31_14), .ow_carry(w_carry_31_14));
wire w_sum_31_12, w_carry_31_12;
math_adder_full FA_31_12(.i_a(w_sum_31_36), .i_b(w_sum_31_34), .i_c(w_sum_31_32), .ow_sum(w_sum_31_12), .ow_carry(w_carry_31_12));
wire w_sum_31_10, w_carry_31_10;
math_adder_full FA_31_10(.i_a(w_sum_31_30), .i_b(w_sum_31_28), .i_c(w_sum_31_26), .ow_sum(w_sum_31_10), .ow_carry(w_carry_31_10));
wire w_sum_31_08, w_carry_31_08;
math_adder_full FA_31_08(.i_a(w_sum_31_24), .i_b(w_sum_31_22), .i_c(w_sum_31_20), .ow_sum(w_sum_31_08), .ow_carry(w_carry_31_08));
wire w_sum_31_06, w_carry_31_06;
math_adder_full FA_31_06(.i_a(w_sum_31_18), .i_b(w_sum_31_16), .i_c(w_sum_31_14), .ow_sum(w_sum_31_06), .ow_carry(w_carry_31_06));
wire w_sum_31_04, w_carry_31_04;
math_adder_full FA_31_04(.i_a(w_sum_31_12), .i_b(w_sum_31_10), .i_c(w_sum_31_08), .ow_sum(w_sum_31_04), .ow_carry(w_carry_31_04));
wire w_sum_31_02, w_carry_31_02;
math_adder_half HA_31_02(.i_a(w_sum_31_06), .i_b(w_sum_31_04), .ow_sum(w_sum_31_02), .ow_carry(w_carry_31_02));
wire w_sum_32_62, w_carry_32_62;
math_adder_full FA_32_62(.i_a(w_pp_01_31), .i_b(w_pp_02_30), .i_c(w_pp_03_29), .ow_sum(w_sum_32_62), .ow_carry(w_carry_32_62));
wire w_sum_32_60, w_carry_32_60;
math_adder_full FA_32_60(.i_a(w_pp_04_28), .i_b(w_pp_05_27), .i_c(w_pp_06_26), .ow_sum(w_sum_32_60), .ow_carry(w_carry_32_60));
wire w_sum_32_58, w_carry_32_58;
math_adder_full FA_32_58(.i_a(w_pp_07_25), .i_b(w_pp_08_24), .i_c(w_pp_09_23), .ow_sum(w_sum_32_58), .ow_carry(w_carry_32_58));
wire w_sum_32_56, w_carry_32_56;
math_adder_full FA_32_56(.i_a(w_pp_10_22), .i_b(w_pp_11_21), .i_c(w_pp_12_20), .ow_sum(w_sum_32_56), .ow_carry(w_carry_32_56));
wire w_sum_32_54, w_carry_32_54;
math_adder_full FA_32_54(.i_a(w_pp_13_19), .i_b(w_pp_14_18), .i_c(w_pp_15_17), .ow_sum(w_sum_32_54), .ow_carry(w_carry_32_54));
wire w_sum_32_52, w_carry_32_52;
math_adder_full FA_32_52(.i_a(w_pp_16_16), .i_b(w_pp_17_15), .i_c(w_pp_18_14), .ow_sum(w_sum_32_52), .ow_carry(w_carry_32_52));
wire w_sum_32_50, w_carry_32_50;
math_adder_full FA_32_50(.i_a(w_pp_19_13), .i_b(w_pp_20_12), .i_c(w_pp_21_11), .ow_sum(w_sum_32_50), .ow_carry(w_carry_32_50));
wire w_sum_32_48, w_carry_32_48;
math_adder_full FA_32_48(.i_a(w_pp_22_10), .i_b(w_pp_23_09), .i_c(w_pp_24_08), .ow_sum(w_sum_32_48), .ow_carry(w_carry_32_48));
wire w_sum_32_46, w_carry_32_46;
math_adder_full FA_32_46(.i_a(w_pp_25_07), .i_b(w_pp_26_06), .i_c(w_pp_27_05), .ow_sum(w_sum_32_46), .ow_carry(w_carry_32_46));
wire w_sum_32_44, w_carry_32_44;
math_adder_full FA_32_44(.i_a(w_pp_28_04), .i_b(w_pp_29_03), .i_c(w_pp_30_02), .ow_sum(w_sum_32_44), .ow_carry(w_carry_32_44));
wire w_sum_32_42, w_carry_32_42;
math_adder_full FA_32_42(.i_a(w_pp_31_01), .i_b(w_carry_31_62), .i_c(w_carry_31_60), .ow_sum(w_sum_32_42), .ow_carry(w_carry_32_42));
wire w_sum_32_40, w_carry_32_40;
math_adder_full FA_32_40(.i_a(w_carry_31_58), .i_b(w_carry_31_56), .i_c(w_carry_31_54), .ow_sum(w_sum_32_40), .ow_carry(w_carry_32_40));
wire w_sum_32_38, w_carry_32_38;
math_adder_full FA_32_38(.i_a(w_carry_31_52), .i_b(w_carry_31_50), .i_c(w_carry_31_48), .ow_sum(w_sum_32_38), .ow_carry(w_carry_32_38));
wire w_sum_32_36, w_carry_32_36;
math_adder_full FA_32_36(.i_a(w_carry_31_46), .i_b(w_carry_31_44), .i_c(w_carry_31_42), .ow_sum(w_sum_32_36), .ow_carry(w_carry_32_36));
wire w_sum_32_34, w_carry_32_34;
math_adder_full FA_32_34(.i_a(w_carry_31_40), .i_b(w_carry_31_38), .i_c(w_carry_31_36), .ow_sum(w_sum_32_34), .ow_carry(w_carry_32_34));
wire w_sum_32_32, w_carry_32_32;
math_adder_full FA_32_32(.i_a(w_carry_31_34), .i_b(w_carry_31_32), .i_c(w_carry_31_30), .ow_sum(w_sum_32_32), .ow_carry(w_carry_32_32));
wire w_sum_32_30, w_carry_32_30;
math_adder_full FA_32_30(.i_a(w_carry_31_28), .i_b(w_carry_31_26), .i_c(w_carry_31_24), .ow_sum(w_sum_32_30), .ow_carry(w_carry_32_30));
wire w_sum_32_28, w_carry_32_28;
math_adder_full FA_32_28(.i_a(w_carry_31_22), .i_b(w_carry_31_20), .i_c(w_carry_31_18), .ow_sum(w_sum_32_28), .ow_carry(w_carry_32_28));
wire w_sum_32_26, w_carry_32_26;
math_adder_full FA_32_26(.i_a(w_carry_31_16), .i_b(w_carry_31_14), .i_c(w_carry_31_12), .ow_sum(w_sum_32_26), .ow_carry(w_carry_32_26));
wire w_sum_32_24, w_carry_32_24;
math_adder_full FA_32_24(.i_a(w_carry_31_10), .i_b(w_carry_31_08), .i_c(w_carry_31_06), .ow_sum(w_sum_32_24), .ow_carry(w_carry_32_24));
wire w_sum_32_22, w_carry_32_22;
math_adder_full FA_32_22(.i_a(w_carry_31_04), .i_b(w_carry_31_02), .i_c(w_sum_32_62), .ow_sum(w_sum_32_22), .ow_carry(w_carry_32_22));
wire w_sum_32_20, w_carry_32_20;
math_adder_full FA_32_20(.i_a(w_sum_32_60), .i_b(w_sum_32_58), .i_c(w_sum_32_56), .ow_sum(w_sum_32_20), .ow_carry(w_carry_32_20));
wire w_sum_32_18, w_carry_32_18;
math_adder_full FA_32_18(.i_a(w_sum_32_54), .i_b(w_sum_32_52), .i_c(w_sum_32_50), .ow_sum(w_sum_32_18), .ow_carry(w_carry_32_18));
wire w_sum_32_16, w_carry_32_16;
math_adder_full FA_32_16(.i_a(w_sum_32_48), .i_b(w_sum_32_46), .i_c(w_sum_32_44), .ow_sum(w_sum_32_16), .ow_carry(w_carry_32_16));
wire w_sum_32_14, w_carry_32_14;
math_adder_full FA_32_14(.i_a(w_sum_32_42), .i_b(w_sum_32_40), .i_c(w_sum_32_38), .ow_sum(w_sum_32_14), .ow_carry(w_carry_32_14));
wire w_sum_32_12, w_carry_32_12;
math_adder_full FA_32_12(.i_a(w_sum_32_36), .i_b(w_sum_32_34), .i_c(w_sum_32_32), .ow_sum(w_sum_32_12), .ow_carry(w_carry_32_12));
wire w_sum_32_10, w_carry_32_10;
math_adder_full FA_32_10(.i_a(w_sum_32_30), .i_b(w_sum_32_28), .i_c(w_sum_32_26), .ow_sum(w_sum_32_10), .ow_carry(w_carry_32_10));
wire w_sum_32_08, w_carry_32_08;
math_adder_full FA_32_08(.i_a(w_sum_32_24), .i_b(w_sum_32_22), .i_c(w_sum_32_20), .ow_sum(w_sum_32_08), .ow_carry(w_carry_32_08));
wire w_sum_32_06, w_carry_32_06;
math_adder_full FA_32_06(.i_a(w_sum_32_18), .i_b(w_sum_32_16), .i_c(w_sum_32_14), .ow_sum(w_sum_32_06), .ow_carry(w_carry_32_06));
wire w_sum_32_04, w_carry_32_04;
math_adder_full FA_32_04(.i_a(w_sum_32_12), .i_b(w_sum_32_10), .i_c(w_sum_32_08), .ow_sum(w_sum_32_04), .ow_carry(w_carry_32_04));
wire w_sum_32_02, w_carry_32_02;
math_adder_half HA_32_02(.i_a(w_sum_32_06), .i_b(w_sum_32_04), .ow_sum(w_sum_32_02), .ow_carry(w_carry_32_02));
wire w_sum_33_61, w_carry_33_61;
math_adder_full FA_33_61(.i_a(w_pp_02_31), .i_b(w_pp_03_30), .i_c(w_pp_04_29), .ow_sum(w_sum_33_61), .ow_carry(w_carry_33_61));
wire w_sum_33_59, w_carry_33_59;
math_adder_full FA_33_59(.i_a(w_pp_05_28), .i_b(w_pp_06_27), .i_c(w_pp_07_26), .ow_sum(w_sum_33_59), .ow_carry(w_carry_33_59));
wire w_sum_33_57, w_carry_33_57;
math_adder_full FA_33_57(.i_a(w_pp_08_25), .i_b(w_pp_09_24), .i_c(w_pp_10_23), .ow_sum(w_sum_33_57), .ow_carry(w_carry_33_57));
wire w_sum_33_55, w_carry_33_55;
math_adder_full FA_33_55(.i_a(w_pp_11_22), .i_b(w_pp_12_21), .i_c(w_pp_13_20), .ow_sum(w_sum_33_55), .ow_carry(w_carry_33_55));
wire w_sum_33_53, w_carry_33_53;
math_adder_full FA_33_53(.i_a(w_pp_14_19), .i_b(w_pp_15_18), .i_c(w_pp_16_17), .ow_sum(w_sum_33_53), .ow_carry(w_carry_33_53));
wire w_sum_33_51, w_carry_33_51;
math_adder_full FA_33_51(.i_a(w_pp_17_16), .i_b(w_pp_18_15), .i_c(w_pp_19_14), .ow_sum(w_sum_33_51), .ow_carry(w_carry_33_51));
wire w_sum_33_49, w_carry_33_49;
math_adder_full FA_33_49(.i_a(w_pp_20_13), .i_b(w_pp_21_12), .i_c(w_pp_22_11), .ow_sum(w_sum_33_49), .ow_carry(w_carry_33_49));
wire w_sum_33_47, w_carry_33_47;
math_adder_full FA_33_47(.i_a(w_pp_23_10), .i_b(w_pp_24_09), .i_c(w_pp_25_08), .ow_sum(w_sum_33_47), .ow_carry(w_carry_33_47));
wire w_sum_33_45, w_carry_33_45;
math_adder_full FA_33_45(.i_a(w_pp_26_07), .i_b(w_pp_27_06), .i_c(w_pp_28_05), .ow_sum(w_sum_33_45), .ow_carry(w_carry_33_45));
wire w_sum_33_43, w_carry_33_43;
math_adder_full FA_33_43(.i_a(w_pp_29_04), .i_b(w_pp_30_03), .i_c(w_pp_31_02), .ow_sum(w_sum_33_43), .ow_carry(w_carry_33_43));
wire w_sum_33_41, w_carry_33_41;
math_adder_full FA_33_41(.i_a(w_carry_32_62), .i_b(w_carry_32_60), .i_c(w_carry_32_58), .ow_sum(w_sum_33_41), .ow_carry(w_carry_33_41));
wire w_sum_33_39, w_carry_33_39;
math_adder_full FA_33_39(.i_a(w_carry_32_56), .i_b(w_carry_32_54), .i_c(w_carry_32_52), .ow_sum(w_sum_33_39), .ow_carry(w_carry_33_39));
wire w_sum_33_37, w_carry_33_37;
math_adder_full FA_33_37(.i_a(w_carry_32_50), .i_b(w_carry_32_48), .i_c(w_carry_32_46), .ow_sum(w_sum_33_37), .ow_carry(w_carry_33_37));
wire w_sum_33_35, w_carry_33_35;
math_adder_full FA_33_35(.i_a(w_carry_32_44), .i_b(w_carry_32_42), .i_c(w_carry_32_40), .ow_sum(w_sum_33_35), .ow_carry(w_carry_33_35));
wire w_sum_33_33, w_carry_33_33;
math_adder_full FA_33_33(.i_a(w_carry_32_38), .i_b(w_carry_32_36), .i_c(w_carry_32_34), .ow_sum(w_sum_33_33), .ow_carry(w_carry_33_33));
wire w_sum_33_31, w_carry_33_31;
math_adder_full FA_33_31(.i_a(w_carry_32_32), .i_b(w_carry_32_30), .i_c(w_carry_32_28), .ow_sum(w_sum_33_31), .ow_carry(w_carry_33_31));
wire w_sum_33_29, w_carry_33_29;
math_adder_full FA_33_29(.i_a(w_carry_32_26), .i_b(w_carry_32_24), .i_c(w_carry_32_22), .ow_sum(w_sum_33_29), .ow_carry(w_carry_33_29));
wire w_sum_33_27, w_carry_33_27;
math_adder_full FA_33_27(.i_a(w_carry_32_20), .i_b(w_carry_32_18), .i_c(w_carry_32_16), .ow_sum(w_sum_33_27), .ow_carry(w_carry_33_27));
wire w_sum_33_25, w_carry_33_25;
math_adder_full FA_33_25(.i_a(w_carry_32_14), .i_b(w_carry_32_12), .i_c(w_carry_32_10), .ow_sum(w_sum_33_25), .ow_carry(w_carry_33_25));
wire w_sum_33_23, w_carry_33_23;
math_adder_full FA_33_23(.i_a(w_carry_32_08), .i_b(w_carry_32_06), .i_c(w_carry_32_04), .ow_sum(w_sum_33_23), .ow_carry(w_carry_33_23));
wire w_sum_33_21, w_carry_33_21;
math_adder_full FA_33_21(.i_a(w_carry_32_02), .i_b(w_sum_33_61), .i_c(w_sum_33_59), .ow_sum(w_sum_33_21), .ow_carry(w_carry_33_21));
wire w_sum_33_19, w_carry_33_19;
math_adder_full FA_33_19(.i_a(w_sum_33_57), .i_b(w_sum_33_55), .i_c(w_sum_33_53), .ow_sum(w_sum_33_19), .ow_carry(w_carry_33_19));
wire w_sum_33_17, w_carry_33_17;
math_adder_full FA_33_17(.i_a(w_sum_33_51), .i_b(w_sum_33_49), .i_c(w_sum_33_47), .ow_sum(w_sum_33_17), .ow_carry(w_carry_33_17));
wire w_sum_33_15, w_carry_33_15;
math_adder_full FA_33_15(.i_a(w_sum_33_45), .i_b(w_sum_33_43), .i_c(w_sum_33_41), .ow_sum(w_sum_33_15), .ow_carry(w_carry_33_15));
wire w_sum_33_13, w_carry_33_13;
math_adder_full FA_33_13(.i_a(w_sum_33_39), .i_b(w_sum_33_37), .i_c(w_sum_33_35), .ow_sum(w_sum_33_13), .ow_carry(w_carry_33_13));
wire w_sum_33_11, w_carry_33_11;
math_adder_full FA_33_11(.i_a(w_sum_33_33), .i_b(w_sum_33_31), .i_c(w_sum_33_29), .ow_sum(w_sum_33_11), .ow_carry(w_carry_33_11));
wire w_sum_33_09, w_carry_33_09;
math_adder_full FA_33_09(.i_a(w_sum_33_27), .i_b(w_sum_33_25), .i_c(w_sum_33_23), .ow_sum(w_sum_33_09), .ow_carry(w_carry_33_09));
wire w_sum_33_07, w_carry_33_07;
math_adder_full FA_33_07(.i_a(w_sum_33_21), .i_b(w_sum_33_19), .i_c(w_sum_33_17), .ow_sum(w_sum_33_07), .ow_carry(w_carry_33_07));
wire w_sum_33_05, w_carry_33_05;
math_adder_full FA_33_05(.i_a(w_sum_33_15), .i_b(w_sum_33_13), .i_c(w_sum_33_11), .ow_sum(w_sum_33_05), .ow_carry(w_carry_33_05));
wire w_sum_33_03, w_carry_33_03;
math_adder_full FA_33_03(.i_a(w_sum_33_09), .i_b(w_sum_33_07), .i_c(w_sum_33_05), .ow_sum(w_sum_33_03), .ow_carry(w_carry_33_03));
wire w_sum_34_59, w_carry_34_59;
math_adder_full FA_34_59(.i_a(w_pp_03_31), .i_b(w_pp_04_30), .i_c(w_pp_05_29), .ow_sum(w_sum_34_59), .ow_carry(w_carry_34_59));
wire w_sum_34_57, w_carry_34_57;
math_adder_full FA_34_57(.i_a(w_pp_06_28), .i_b(w_pp_07_27), .i_c(w_pp_08_26), .ow_sum(w_sum_34_57), .ow_carry(w_carry_34_57));
wire w_sum_34_55, w_carry_34_55;
math_adder_full FA_34_55(.i_a(w_pp_09_25), .i_b(w_pp_10_24), .i_c(w_pp_11_23), .ow_sum(w_sum_34_55), .ow_carry(w_carry_34_55));
wire w_sum_34_53, w_carry_34_53;
math_adder_full FA_34_53(.i_a(w_pp_12_22), .i_b(w_pp_13_21), .i_c(w_pp_14_20), .ow_sum(w_sum_34_53), .ow_carry(w_carry_34_53));
wire w_sum_34_51, w_carry_34_51;
math_adder_full FA_34_51(.i_a(w_pp_15_19), .i_b(w_pp_16_18), .i_c(w_pp_17_17), .ow_sum(w_sum_34_51), .ow_carry(w_carry_34_51));
wire w_sum_34_49, w_carry_34_49;
math_adder_full FA_34_49(.i_a(w_pp_18_16), .i_b(w_pp_19_15), .i_c(w_pp_20_14), .ow_sum(w_sum_34_49), .ow_carry(w_carry_34_49));
wire w_sum_34_47, w_carry_34_47;
math_adder_full FA_34_47(.i_a(w_pp_21_13), .i_b(w_pp_22_12), .i_c(w_pp_23_11), .ow_sum(w_sum_34_47), .ow_carry(w_carry_34_47));
wire w_sum_34_45, w_carry_34_45;
math_adder_full FA_34_45(.i_a(w_pp_24_10), .i_b(w_pp_25_09), .i_c(w_pp_26_08), .ow_sum(w_sum_34_45), .ow_carry(w_carry_34_45));
wire w_sum_34_43, w_carry_34_43;
math_adder_full FA_34_43(.i_a(w_pp_27_07), .i_b(w_pp_28_06), .i_c(w_pp_29_05), .ow_sum(w_sum_34_43), .ow_carry(w_carry_34_43));
wire w_sum_34_41, w_carry_34_41;
math_adder_full FA_34_41(.i_a(w_pp_30_04), .i_b(w_pp_31_03), .i_c(w_carry_33_61), .ow_sum(w_sum_34_41), .ow_carry(w_carry_34_41));
wire w_sum_34_39, w_carry_34_39;
math_adder_full FA_34_39(.i_a(w_carry_33_59), .i_b(w_carry_33_57), .i_c(w_carry_33_55), .ow_sum(w_sum_34_39), .ow_carry(w_carry_34_39));
wire w_sum_34_37, w_carry_34_37;
math_adder_full FA_34_37(.i_a(w_carry_33_53), .i_b(w_carry_33_51), .i_c(w_carry_33_49), .ow_sum(w_sum_34_37), .ow_carry(w_carry_34_37));
wire w_sum_34_35, w_carry_34_35;
math_adder_full FA_34_35(.i_a(w_carry_33_47), .i_b(w_carry_33_45), .i_c(w_carry_33_43), .ow_sum(w_sum_34_35), .ow_carry(w_carry_34_35));
wire w_sum_34_33, w_carry_34_33;
math_adder_full FA_34_33(.i_a(w_carry_33_41), .i_b(w_carry_33_39), .i_c(w_carry_33_37), .ow_sum(w_sum_34_33), .ow_carry(w_carry_34_33));
wire w_sum_34_31, w_carry_34_31;
math_adder_full FA_34_31(.i_a(w_carry_33_35), .i_b(w_carry_33_33), .i_c(w_carry_33_31), .ow_sum(w_sum_34_31), .ow_carry(w_carry_34_31));
wire w_sum_34_29, w_carry_34_29;
math_adder_full FA_34_29(.i_a(w_carry_33_29), .i_b(w_carry_33_27), .i_c(w_carry_33_25), .ow_sum(w_sum_34_29), .ow_carry(w_carry_34_29));
wire w_sum_34_27, w_carry_34_27;
math_adder_full FA_34_27(.i_a(w_carry_33_23), .i_b(w_carry_33_21), .i_c(w_carry_33_19), .ow_sum(w_sum_34_27), .ow_carry(w_carry_34_27));
wire w_sum_34_25, w_carry_34_25;
math_adder_full FA_34_25(.i_a(w_carry_33_17), .i_b(w_carry_33_15), .i_c(w_carry_33_13), .ow_sum(w_sum_34_25), .ow_carry(w_carry_34_25));
wire w_sum_34_23, w_carry_34_23;
math_adder_full FA_34_23(.i_a(w_carry_33_11), .i_b(w_carry_33_09), .i_c(w_carry_33_07), .ow_sum(w_sum_34_23), .ow_carry(w_carry_34_23));
wire w_sum_34_21, w_carry_34_21;
math_adder_full FA_34_21(.i_a(w_carry_33_05), .i_b(w_carry_33_03), .i_c(w_sum_34_59), .ow_sum(w_sum_34_21), .ow_carry(w_carry_34_21));
wire w_sum_34_19, w_carry_34_19;
math_adder_full FA_34_19(.i_a(w_sum_34_57), .i_b(w_sum_34_55), .i_c(w_sum_34_53), .ow_sum(w_sum_34_19), .ow_carry(w_carry_34_19));
wire w_sum_34_17, w_carry_34_17;
math_adder_full FA_34_17(.i_a(w_sum_34_51), .i_b(w_sum_34_49), .i_c(w_sum_34_47), .ow_sum(w_sum_34_17), .ow_carry(w_carry_34_17));
wire w_sum_34_15, w_carry_34_15;
math_adder_full FA_34_15(.i_a(w_sum_34_45), .i_b(w_sum_34_43), .i_c(w_sum_34_41), .ow_sum(w_sum_34_15), .ow_carry(w_carry_34_15));
wire w_sum_34_13, w_carry_34_13;
math_adder_full FA_34_13(.i_a(w_sum_34_39), .i_b(w_sum_34_37), .i_c(w_sum_34_35), .ow_sum(w_sum_34_13), .ow_carry(w_carry_34_13));
wire w_sum_34_11, w_carry_34_11;
math_adder_full FA_34_11(.i_a(w_sum_34_33), .i_b(w_sum_34_31), .i_c(w_sum_34_29), .ow_sum(w_sum_34_11), .ow_carry(w_carry_34_11));
wire w_sum_34_09, w_carry_34_09;
math_adder_full FA_34_09(.i_a(w_sum_34_27), .i_b(w_sum_34_25), .i_c(w_sum_34_23), .ow_sum(w_sum_34_09), .ow_carry(w_carry_34_09));
wire w_sum_34_07, w_carry_34_07;
math_adder_full FA_34_07(.i_a(w_sum_34_21), .i_b(w_sum_34_19), .i_c(w_sum_34_17), .ow_sum(w_sum_34_07), .ow_carry(w_carry_34_07));
wire w_sum_34_05, w_carry_34_05;
math_adder_full FA_34_05(.i_a(w_sum_34_15), .i_b(w_sum_34_13), .i_c(w_sum_34_11), .ow_sum(w_sum_34_05), .ow_carry(w_carry_34_05));
wire w_sum_34_03, w_carry_34_03;
math_adder_full FA_34_03(.i_a(w_sum_34_09), .i_b(w_sum_34_07), .i_c(w_sum_34_05), .ow_sum(w_sum_34_03), .ow_carry(w_carry_34_03));
wire w_sum_35_57, w_carry_35_57;
math_adder_full FA_35_57(.i_a(w_pp_04_31), .i_b(w_pp_05_30), .i_c(w_pp_06_29), .ow_sum(w_sum_35_57), .ow_carry(w_carry_35_57));
wire w_sum_35_55, w_carry_35_55;
math_adder_full FA_35_55(.i_a(w_pp_07_28), .i_b(w_pp_08_27), .i_c(w_pp_09_26), .ow_sum(w_sum_35_55), .ow_carry(w_carry_35_55));
wire w_sum_35_53, w_carry_35_53;
math_adder_full FA_35_53(.i_a(w_pp_10_25), .i_b(w_pp_11_24), .i_c(w_pp_12_23), .ow_sum(w_sum_35_53), .ow_carry(w_carry_35_53));
wire w_sum_35_51, w_carry_35_51;
math_adder_full FA_35_51(.i_a(w_pp_13_22), .i_b(w_pp_14_21), .i_c(w_pp_15_20), .ow_sum(w_sum_35_51), .ow_carry(w_carry_35_51));
wire w_sum_35_49, w_carry_35_49;
math_adder_full FA_35_49(.i_a(w_pp_16_19), .i_b(w_pp_17_18), .i_c(w_pp_18_17), .ow_sum(w_sum_35_49), .ow_carry(w_carry_35_49));
wire w_sum_35_47, w_carry_35_47;
math_adder_full FA_35_47(.i_a(w_pp_19_16), .i_b(w_pp_20_15), .i_c(w_pp_21_14), .ow_sum(w_sum_35_47), .ow_carry(w_carry_35_47));
wire w_sum_35_45, w_carry_35_45;
math_adder_full FA_35_45(.i_a(w_pp_22_13), .i_b(w_pp_23_12), .i_c(w_pp_24_11), .ow_sum(w_sum_35_45), .ow_carry(w_carry_35_45));
wire w_sum_35_43, w_carry_35_43;
math_adder_full FA_35_43(.i_a(w_pp_25_10), .i_b(w_pp_26_09), .i_c(w_pp_27_08), .ow_sum(w_sum_35_43), .ow_carry(w_carry_35_43));
wire w_sum_35_41, w_carry_35_41;
math_adder_full FA_35_41(.i_a(w_pp_28_07), .i_b(w_pp_29_06), .i_c(w_pp_30_05), .ow_sum(w_sum_35_41), .ow_carry(w_carry_35_41));
wire w_sum_35_39, w_carry_35_39;
math_adder_full FA_35_39(.i_a(w_pp_31_04), .i_b(w_carry_34_59), .i_c(w_carry_34_57), .ow_sum(w_sum_35_39), .ow_carry(w_carry_35_39));
wire w_sum_35_37, w_carry_35_37;
math_adder_full FA_35_37(.i_a(w_carry_34_55), .i_b(w_carry_34_53), .i_c(w_carry_34_51), .ow_sum(w_sum_35_37), .ow_carry(w_carry_35_37));
wire w_sum_35_35, w_carry_35_35;
math_adder_full FA_35_35(.i_a(w_carry_34_49), .i_b(w_carry_34_47), .i_c(w_carry_34_45), .ow_sum(w_sum_35_35), .ow_carry(w_carry_35_35));
wire w_sum_35_33, w_carry_35_33;
math_adder_full FA_35_33(.i_a(w_carry_34_43), .i_b(w_carry_34_41), .i_c(w_carry_34_39), .ow_sum(w_sum_35_33), .ow_carry(w_carry_35_33));
wire w_sum_35_31, w_carry_35_31;
math_adder_full FA_35_31(.i_a(w_carry_34_37), .i_b(w_carry_34_35), .i_c(w_carry_34_33), .ow_sum(w_sum_35_31), .ow_carry(w_carry_35_31));
wire w_sum_35_29, w_carry_35_29;
math_adder_full FA_35_29(.i_a(w_carry_34_31), .i_b(w_carry_34_29), .i_c(w_carry_34_27), .ow_sum(w_sum_35_29), .ow_carry(w_carry_35_29));
wire w_sum_35_27, w_carry_35_27;
math_adder_full FA_35_27(.i_a(w_carry_34_25), .i_b(w_carry_34_23), .i_c(w_carry_34_21), .ow_sum(w_sum_35_27), .ow_carry(w_carry_35_27));
wire w_sum_35_25, w_carry_35_25;
math_adder_full FA_35_25(.i_a(w_carry_34_19), .i_b(w_carry_34_17), .i_c(w_carry_34_15), .ow_sum(w_sum_35_25), .ow_carry(w_carry_35_25));
wire w_sum_35_23, w_carry_35_23;
math_adder_full FA_35_23(.i_a(w_carry_34_13), .i_b(w_carry_34_11), .i_c(w_carry_34_09), .ow_sum(w_sum_35_23), .ow_carry(w_carry_35_23));
wire w_sum_35_21, w_carry_35_21;
math_adder_full FA_35_21(.i_a(w_carry_34_07), .i_b(w_carry_34_05), .i_c(w_carry_34_03), .ow_sum(w_sum_35_21), .ow_carry(w_carry_35_21));
wire w_sum_35_19, w_carry_35_19;
math_adder_full FA_35_19(.i_a(w_sum_35_57), .i_b(w_sum_35_55), .i_c(w_sum_35_53), .ow_sum(w_sum_35_19), .ow_carry(w_carry_35_19));
wire w_sum_35_17, w_carry_35_17;
math_adder_full FA_35_17(.i_a(w_sum_35_51), .i_b(w_sum_35_49), .i_c(w_sum_35_47), .ow_sum(w_sum_35_17), .ow_carry(w_carry_35_17));
wire w_sum_35_15, w_carry_35_15;
math_adder_full FA_35_15(.i_a(w_sum_35_45), .i_b(w_sum_35_43), .i_c(w_sum_35_41), .ow_sum(w_sum_35_15), .ow_carry(w_carry_35_15));
wire w_sum_35_13, w_carry_35_13;
math_adder_full FA_35_13(.i_a(w_sum_35_39), .i_b(w_sum_35_37), .i_c(w_sum_35_35), .ow_sum(w_sum_35_13), .ow_carry(w_carry_35_13));
wire w_sum_35_11, w_carry_35_11;
math_adder_full FA_35_11(.i_a(w_sum_35_33), .i_b(w_sum_35_31), .i_c(w_sum_35_29), .ow_sum(w_sum_35_11), .ow_carry(w_carry_35_11));
wire w_sum_35_09, w_carry_35_09;
math_adder_full FA_35_09(.i_a(w_sum_35_27), .i_b(w_sum_35_25), .i_c(w_sum_35_23), .ow_sum(w_sum_35_09), .ow_carry(w_carry_35_09));
wire w_sum_35_07, w_carry_35_07;
math_adder_full FA_35_07(.i_a(w_sum_35_21), .i_b(w_sum_35_19), .i_c(w_sum_35_17), .ow_sum(w_sum_35_07), .ow_carry(w_carry_35_07));
wire w_sum_35_05, w_carry_35_05;
math_adder_full FA_35_05(.i_a(w_sum_35_15), .i_b(w_sum_35_13), .i_c(w_sum_35_11), .ow_sum(w_sum_35_05), .ow_carry(w_carry_35_05));
wire w_sum_35_03, w_carry_35_03;
math_adder_full FA_35_03(.i_a(w_sum_35_09), .i_b(w_sum_35_07), .i_c(w_sum_35_05), .ow_sum(w_sum_35_03), .ow_carry(w_carry_35_03));
wire w_sum_36_55, w_carry_36_55;
math_adder_full FA_36_55(.i_a(w_pp_05_31), .i_b(w_pp_06_30), .i_c(w_pp_07_29), .ow_sum(w_sum_36_55), .ow_carry(w_carry_36_55));
wire w_sum_36_53, w_carry_36_53;
math_adder_full FA_36_53(.i_a(w_pp_08_28), .i_b(w_pp_09_27), .i_c(w_pp_10_26), .ow_sum(w_sum_36_53), .ow_carry(w_carry_36_53));
wire w_sum_36_51, w_carry_36_51;
math_adder_full FA_36_51(.i_a(w_pp_11_25), .i_b(w_pp_12_24), .i_c(w_pp_13_23), .ow_sum(w_sum_36_51), .ow_carry(w_carry_36_51));
wire w_sum_36_49, w_carry_36_49;
math_adder_full FA_36_49(.i_a(w_pp_14_22), .i_b(w_pp_15_21), .i_c(w_pp_16_20), .ow_sum(w_sum_36_49), .ow_carry(w_carry_36_49));
wire w_sum_36_47, w_carry_36_47;
math_adder_full FA_36_47(.i_a(w_pp_17_19), .i_b(w_pp_18_18), .i_c(w_pp_19_17), .ow_sum(w_sum_36_47), .ow_carry(w_carry_36_47));
wire w_sum_36_45, w_carry_36_45;
math_adder_full FA_36_45(.i_a(w_pp_20_16), .i_b(w_pp_21_15), .i_c(w_pp_22_14), .ow_sum(w_sum_36_45), .ow_carry(w_carry_36_45));
wire w_sum_36_43, w_carry_36_43;
math_adder_full FA_36_43(.i_a(w_pp_23_13), .i_b(w_pp_24_12), .i_c(w_pp_25_11), .ow_sum(w_sum_36_43), .ow_carry(w_carry_36_43));
wire w_sum_36_41, w_carry_36_41;
math_adder_full FA_36_41(.i_a(w_pp_26_10), .i_b(w_pp_27_09), .i_c(w_pp_28_08), .ow_sum(w_sum_36_41), .ow_carry(w_carry_36_41));
wire w_sum_36_39, w_carry_36_39;
math_adder_full FA_36_39(.i_a(w_pp_29_07), .i_b(w_pp_30_06), .i_c(w_pp_31_05), .ow_sum(w_sum_36_39), .ow_carry(w_carry_36_39));
wire w_sum_36_37, w_carry_36_37;
math_adder_full FA_36_37(.i_a(w_carry_35_57), .i_b(w_carry_35_55), .i_c(w_carry_35_53), .ow_sum(w_sum_36_37), .ow_carry(w_carry_36_37));
wire w_sum_36_35, w_carry_36_35;
math_adder_full FA_36_35(.i_a(w_carry_35_51), .i_b(w_carry_35_49), .i_c(w_carry_35_47), .ow_sum(w_sum_36_35), .ow_carry(w_carry_36_35));
wire w_sum_36_33, w_carry_36_33;
math_adder_full FA_36_33(.i_a(w_carry_35_45), .i_b(w_carry_35_43), .i_c(w_carry_35_41), .ow_sum(w_sum_36_33), .ow_carry(w_carry_36_33));
wire w_sum_36_31, w_carry_36_31;
math_adder_full FA_36_31(.i_a(w_carry_35_39), .i_b(w_carry_35_37), .i_c(w_carry_35_35), .ow_sum(w_sum_36_31), .ow_carry(w_carry_36_31));
wire w_sum_36_29, w_carry_36_29;
math_adder_full FA_36_29(.i_a(w_carry_35_33), .i_b(w_carry_35_31), .i_c(w_carry_35_29), .ow_sum(w_sum_36_29), .ow_carry(w_carry_36_29));
wire w_sum_36_27, w_carry_36_27;
math_adder_full FA_36_27(.i_a(w_carry_35_27), .i_b(w_carry_35_25), .i_c(w_carry_35_23), .ow_sum(w_sum_36_27), .ow_carry(w_carry_36_27));
wire w_sum_36_25, w_carry_36_25;
math_adder_full FA_36_25(.i_a(w_carry_35_21), .i_b(w_carry_35_19), .i_c(w_carry_35_17), .ow_sum(w_sum_36_25), .ow_carry(w_carry_36_25));
wire w_sum_36_23, w_carry_36_23;
math_adder_full FA_36_23(.i_a(w_carry_35_15), .i_b(w_carry_35_13), .i_c(w_carry_35_11), .ow_sum(w_sum_36_23), .ow_carry(w_carry_36_23));
wire w_sum_36_21, w_carry_36_21;
math_adder_full FA_36_21(.i_a(w_carry_35_09), .i_b(w_carry_35_07), .i_c(w_carry_35_05), .ow_sum(w_sum_36_21), .ow_carry(w_carry_36_21));
wire w_sum_36_19, w_carry_36_19;
math_adder_full FA_36_19(.i_a(w_carry_35_03), .i_b(w_sum_36_55), .i_c(w_sum_36_53), .ow_sum(w_sum_36_19), .ow_carry(w_carry_36_19));
wire w_sum_36_17, w_carry_36_17;
math_adder_full FA_36_17(.i_a(w_sum_36_51), .i_b(w_sum_36_49), .i_c(w_sum_36_47), .ow_sum(w_sum_36_17), .ow_carry(w_carry_36_17));
wire w_sum_36_15, w_carry_36_15;
math_adder_full FA_36_15(.i_a(w_sum_36_45), .i_b(w_sum_36_43), .i_c(w_sum_36_41), .ow_sum(w_sum_36_15), .ow_carry(w_carry_36_15));
wire w_sum_36_13, w_carry_36_13;
math_adder_full FA_36_13(.i_a(w_sum_36_39), .i_b(w_sum_36_37), .i_c(w_sum_36_35), .ow_sum(w_sum_36_13), .ow_carry(w_carry_36_13));
wire w_sum_36_11, w_carry_36_11;
math_adder_full FA_36_11(.i_a(w_sum_36_33), .i_b(w_sum_36_31), .i_c(w_sum_36_29), .ow_sum(w_sum_36_11), .ow_carry(w_carry_36_11));
wire w_sum_36_09, w_carry_36_09;
math_adder_full FA_36_09(.i_a(w_sum_36_27), .i_b(w_sum_36_25), .i_c(w_sum_36_23), .ow_sum(w_sum_36_09), .ow_carry(w_carry_36_09));
wire w_sum_36_07, w_carry_36_07;
math_adder_full FA_36_07(.i_a(w_sum_36_21), .i_b(w_sum_36_19), .i_c(w_sum_36_17), .ow_sum(w_sum_36_07), .ow_carry(w_carry_36_07));
wire w_sum_36_05, w_carry_36_05;
math_adder_full FA_36_05(.i_a(w_sum_36_15), .i_b(w_sum_36_13), .i_c(w_sum_36_11), .ow_sum(w_sum_36_05), .ow_carry(w_carry_36_05));
wire w_sum_36_03, w_carry_36_03;
math_adder_full FA_36_03(.i_a(w_sum_36_09), .i_b(w_sum_36_07), .i_c(w_sum_36_05), .ow_sum(w_sum_36_03), .ow_carry(w_carry_36_03));
wire w_sum_37_53, w_carry_37_53;
math_adder_full FA_37_53(.i_a(w_pp_06_31), .i_b(w_pp_07_30), .i_c(w_pp_08_29), .ow_sum(w_sum_37_53), .ow_carry(w_carry_37_53));
wire w_sum_37_51, w_carry_37_51;
math_adder_full FA_37_51(.i_a(w_pp_09_28), .i_b(w_pp_10_27), .i_c(w_pp_11_26), .ow_sum(w_sum_37_51), .ow_carry(w_carry_37_51));
wire w_sum_37_49, w_carry_37_49;
math_adder_full FA_37_49(.i_a(w_pp_12_25), .i_b(w_pp_13_24), .i_c(w_pp_14_23), .ow_sum(w_sum_37_49), .ow_carry(w_carry_37_49));
wire w_sum_37_47, w_carry_37_47;
math_adder_full FA_37_47(.i_a(w_pp_15_22), .i_b(w_pp_16_21), .i_c(w_pp_17_20), .ow_sum(w_sum_37_47), .ow_carry(w_carry_37_47));
wire w_sum_37_45, w_carry_37_45;
math_adder_full FA_37_45(.i_a(w_pp_18_19), .i_b(w_pp_19_18), .i_c(w_pp_20_17), .ow_sum(w_sum_37_45), .ow_carry(w_carry_37_45));
wire w_sum_37_43, w_carry_37_43;
math_adder_full FA_37_43(.i_a(w_pp_21_16), .i_b(w_pp_22_15), .i_c(w_pp_23_14), .ow_sum(w_sum_37_43), .ow_carry(w_carry_37_43));
wire w_sum_37_41, w_carry_37_41;
math_adder_full FA_37_41(.i_a(w_pp_24_13), .i_b(w_pp_25_12), .i_c(w_pp_26_11), .ow_sum(w_sum_37_41), .ow_carry(w_carry_37_41));
wire w_sum_37_39, w_carry_37_39;
math_adder_full FA_37_39(.i_a(w_pp_27_10), .i_b(w_pp_28_09), .i_c(w_pp_29_08), .ow_sum(w_sum_37_39), .ow_carry(w_carry_37_39));
wire w_sum_37_37, w_carry_37_37;
math_adder_full FA_37_37(.i_a(w_pp_30_07), .i_b(w_pp_31_06), .i_c(w_carry_36_55), .ow_sum(w_sum_37_37), .ow_carry(w_carry_37_37));
wire w_sum_37_35, w_carry_37_35;
math_adder_full FA_37_35(.i_a(w_carry_36_53), .i_b(w_carry_36_51), .i_c(w_carry_36_49), .ow_sum(w_sum_37_35), .ow_carry(w_carry_37_35));
wire w_sum_37_33, w_carry_37_33;
math_adder_full FA_37_33(.i_a(w_carry_36_47), .i_b(w_carry_36_45), .i_c(w_carry_36_43), .ow_sum(w_sum_37_33), .ow_carry(w_carry_37_33));
wire w_sum_37_31, w_carry_37_31;
math_adder_full FA_37_31(.i_a(w_carry_36_41), .i_b(w_carry_36_39), .i_c(w_carry_36_37), .ow_sum(w_sum_37_31), .ow_carry(w_carry_37_31));
wire w_sum_37_29, w_carry_37_29;
math_adder_full FA_37_29(.i_a(w_carry_36_35), .i_b(w_carry_36_33), .i_c(w_carry_36_31), .ow_sum(w_sum_37_29), .ow_carry(w_carry_37_29));
wire w_sum_37_27, w_carry_37_27;
math_adder_full FA_37_27(.i_a(w_carry_36_29), .i_b(w_carry_36_27), .i_c(w_carry_36_25), .ow_sum(w_sum_37_27), .ow_carry(w_carry_37_27));
wire w_sum_37_25, w_carry_37_25;
math_adder_full FA_37_25(.i_a(w_carry_36_23), .i_b(w_carry_36_21), .i_c(w_carry_36_19), .ow_sum(w_sum_37_25), .ow_carry(w_carry_37_25));
wire w_sum_37_23, w_carry_37_23;
math_adder_full FA_37_23(.i_a(w_carry_36_17), .i_b(w_carry_36_15), .i_c(w_carry_36_13), .ow_sum(w_sum_37_23), .ow_carry(w_carry_37_23));
wire w_sum_37_21, w_carry_37_21;
math_adder_full FA_37_21(.i_a(w_carry_36_11), .i_b(w_carry_36_09), .i_c(w_carry_36_07), .ow_sum(w_sum_37_21), .ow_carry(w_carry_37_21));
wire w_sum_37_19, w_carry_37_19;
math_adder_full FA_37_19(.i_a(w_carry_36_05), .i_b(w_carry_36_03), .i_c(w_sum_37_53), .ow_sum(w_sum_37_19), .ow_carry(w_carry_37_19));
wire w_sum_37_17, w_carry_37_17;
math_adder_full FA_37_17(.i_a(w_sum_37_51), .i_b(w_sum_37_49), .i_c(w_sum_37_47), .ow_sum(w_sum_37_17), .ow_carry(w_carry_37_17));
wire w_sum_37_15, w_carry_37_15;
math_adder_full FA_37_15(.i_a(w_sum_37_45), .i_b(w_sum_37_43), .i_c(w_sum_37_41), .ow_sum(w_sum_37_15), .ow_carry(w_carry_37_15));
wire w_sum_37_13, w_carry_37_13;
math_adder_full FA_37_13(.i_a(w_sum_37_39), .i_b(w_sum_37_37), .i_c(w_sum_37_35), .ow_sum(w_sum_37_13), .ow_carry(w_carry_37_13));
wire w_sum_37_11, w_carry_37_11;
math_adder_full FA_37_11(.i_a(w_sum_37_33), .i_b(w_sum_37_31), .i_c(w_sum_37_29), .ow_sum(w_sum_37_11), .ow_carry(w_carry_37_11));
wire w_sum_37_09, w_carry_37_09;
math_adder_full FA_37_09(.i_a(w_sum_37_27), .i_b(w_sum_37_25), .i_c(w_sum_37_23), .ow_sum(w_sum_37_09), .ow_carry(w_carry_37_09));
wire w_sum_37_07, w_carry_37_07;
math_adder_full FA_37_07(.i_a(w_sum_37_21), .i_b(w_sum_37_19), .i_c(w_sum_37_17), .ow_sum(w_sum_37_07), .ow_carry(w_carry_37_07));
wire w_sum_37_05, w_carry_37_05;
math_adder_full FA_37_05(.i_a(w_sum_37_15), .i_b(w_sum_37_13), .i_c(w_sum_37_11), .ow_sum(w_sum_37_05), .ow_carry(w_carry_37_05));
wire w_sum_37_03, w_carry_37_03;
math_adder_full FA_37_03(.i_a(w_sum_37_09), .i_b(w_sum_37_07), .i_c(w_sum_37_05), .ow_sum(w_sum_37_03), .ow_carry(w_carry_37_03));
wire w_sum_38_51, w_carry_38_51;
math_adder_full FA_38_51(.i_a(w_pp_07_31), .i_b(w_pp_08_30), .i_c(w_pp_09_29), .ow_sum(w_sum_38_51), .ow_carry(w_carry_38_51));
wire w_sum_38_49, w_carry_38_49;
math_adder_full FA_38_49(.i_a(w_pp_10_28), .i_b(w_pp_11_27), .i_c(w_pp_12_26), .ow_sum(w_sum_38_49), .ow_carry(w_carry_38_49));
wire w_sum_38_47, w_carry_38_47;
math_adder_full FA_38_47(.i_a(w_pp_13_25), .i_b(w_pp_14_24), .i_c(w_pp_15_23), .ow_sum(w_sum_38_47), .ow_carry(w_carry_38_47));
wire w_sum_38_45, w_carry_38_45;
math_adder_full FA_38_45(.i_a(w_pp_16_22), .i_b(w_pp_17_21), .i_c(w_pp_18_20), .ow_sum(w_sum_38_45), .ow_carry(w_carry_38_45));
wire w_sum_38_43, w_carry_38_43;
math_adder_full FA_38_43(.i_a(w_pp_19_19), .i_b(w_pp_20_18), .i_c(w_pp_21_17), .ow_sum(w_sum_38_43), .ow_carry(w_carry_38_43));
wire w_sum_38_41, w_carry_38_41;
math_adder_full FA_38_41(.i_a(w_pp_22_16), .i_b(w_pp_23_15), .i_c(w_pp_24_14), .ow_sum(w_sum_38_41), .ow_carry(w_carry_38_41));
wire w_sum_38_39, w_carry_38_39;
math_adder_full FA_38_39(.i_a(w_pp_25_13), .i_b(w_pp_26_12), .i_c(w_pp_27_11), .ow_sum(w_sum_38_39), .ow_carry(w_carry_38_39));
wire w_sum_38_37, w_carry_38_37;
math_adder_full FA_38_37(.i_a(w_pp_28_10), .i_b(w_pp_29_09), .i_c(w_pp_30_08), .ow_sum(w_sum_38_37), .ow_carry(w_carry_38_37));
wire w_sum_38_35, w_carry_38_35;
math_adder_full FA_38_35(.i_a(w_pp_31_07), .i_b(w_carry_37_53), .i_c(w_carry_37_51), .ow_sum(w_sum_38_35), .ow_carry(w_carry_38_35));
wire w_sum_38_33, w_carry_38_33;
math_adder_full FA_38_33(.i_a(w_carry_37_49), .i_b(w_carry_37_47), .i_c(w_carry_37_45), .ow_sum(w_sum_38_33), .ow_carry(w_carry_38_33));
wire w_sum_38_31, w_carry_38_31;
math_adder_full FA_38_31(.i_a(w_carry_37_43), .i_b(w_carry_37_41), .i_c(w_carry_37_39), .ow_sum(w_sum_38_31), .ow_carry(w_carry_38_31));
wire w_sum_38_29, w_carry_38_29;
math_adder_full FA_38_29(.i_a(w_carry_37_37), .i_b(w_carry_37_35), .i_c(w_carry_37_33), .ow_sum(w_sum_38_29), .ow_carry(w_carry_38_29));
wire w_sum_38_27, w_carry_38_27;
math_adder_full FA_38_27(.i_a(w_carry_37_31), .i_b(w_carry_37_29), .i_c(w_carry_37_27), .ow_sum(w_sum_38_27), .ow_carry(w_carry_38_27));
wire w_sum_38_25, w_carry_38_25;
math_adder_full FA_38_25(.i_a(w_carry_37_25), .i_b(w_carry_37_23), .i_c(w_carry_37_21), .ow_sum(w_sum_38_25), .ow_carry(w_carry_38_25));
wire w_sum_38_23, w_carry_38_23;
math_adder_full FA_38_23(.i_a(w_carry_37_19), .i_b(w_carry_37_17), .i_c(w_carry_37_15), .ow_sum(w_sum_38_23), .ow_carry(w_carry_38_23));
wire w_sum_38_21, w_carry_38_21;
math_adder_full FA_38_21(.i_a(w_carry_37_13), .i_b(w_carry_37_11), .i_c(w_carry_37_09), .ow_sum(w_sum_38_21), .ow_carry(w_carry_38_21));
wire w_sum_38_19, w_carry_38_19;
math_adder_full FA_38_19(.i_a(w_carry_37_07), .i_b(w_carry_37_05), .i_c(w_carry_37_03), .ow_sum(w_sum_38_19), .ow_carry(w_carry_38_19));
wire w_sum_38_17, w_carry_38_17;
math_adder_full FA_38_17(.i_a(w_sum_38_51), .i_b(w_sum_38_49), .i_c(w_sum_38_47), .ow_sum(w_sum_38_17), .ow_carry(w_carry_38_17));
wire w_sum_38_15, w_carry_38_15;
math_adder_full FA_38_15(.i_a(w_sum_38_45), .i_b(w_sum_38_43), .i_c(w_sum_38_41), .ow_sum(w_sum_38_15), .ow_carry(w_carry_38_15));
wire w_sum_38_13, w_carry_38_13;
math_adder_full FA_38_13(.i_a(w_sum_38_39), .i_b(w_sum_38_37), .i_c(w_sum_38_35), .ow_sum(w_sum_38_13), .ow_carry(w_carry_38_13));
wire w_sum_38_11, w_carry_38_11;
math_adder_full FA_38_11(.i_a(w_sum_38_33), .i_b(w_sum_38_31), .i_c(w_sum_38_29), .ow_sum(w_sum_38_11), .ow_carry(w_carry_38_11));
wire w_sum_38_09, w_carry_38_09;
math_adder_full FA_38_09(.i_a(w_sum_38_27), .i_b(w_sum_38_25), .i_c(w_sum_38_23), .ow_sum(w_sum_38_09), .ow_carry(w_carry_38_09));
wire w_sum_38_07, w_carry_38_07;
math_adder_full FA_38_07(.i_a(w_sum_38_21), .i_b(w_sum_38_19), .i_c(w_sum_38_17), .ow_sum(w_sum_38_07), .ow_carry(w_carry_38_07));
wire w_sum_38_05, w_carry_38_05;
math_adder_full FA_38_05(.i_a(w_sum_38_15), .i_b(w_sum_38_13), .i_c(w_sum_38_11), .ow_sum(w_sum_38_05), .ow_carry(w_carry_38_05));
wire w_sum_38_03, w_carry_38_03;
math_adder_full FA_38_03(.i_a(w_sum_38_09), .i_b(w_sum_38_07), .i_c(w_sum_38_05), .ow_sum(w_sum_38_03), .ow_carry(w_carry_38_03));
wire w_sum_39_49, w_carry_39_49;
math_adder_full FA_39_49(.i_a(w_pp_08_31), .i_b(w_pp_09_30), .i_c(w_pp_10_29), .ow_sum(w_sum_39_49), .ow_carry(w_carry_39_49));
wire w_sum_39_47, w_carry_39_47;
math_adder_full FA_39_47(.i_a(w_pp_11_28), .i_b(w_pp_12_27), .i_c(w_pp_13_26), .ow_sum(w_sum_39_47), .ow_carry(w_carry_39_47));
wire w_sum_39_45, w_carry_39_45;
math_adder_full FA_39_45(.i_a(w_pp_14_25), .i_b(w_pp_15_24), .i_c(w_pp_16_23), .ow_sum(w_sum_39_45), .ow_carry(w_carry_39_45));
wire w_sum_39_43, w_carry_39_43;
math_adder_full FA_39_43(.i_a(w_pp_17_22), .i_b(w_pp_18_21), .i_c(w_pp_19_20), .ow_sum(w_sum_39_43), .ow_carry(w_carry_39_43));
wire w_sum_39_41, w_carry_39_41;
math_adder_full FA_39_41(.i_a(w_pp_20_19), .i_b(w_pp_21_18), .i_c(w_pp_22_17), .ow_sum(w_sum_39_41), .ow_carry(w_carry_39_41));
wire w_sum_39_39, w_carry_39_39;
math_adder_full FA_39_39(.i_a(w_pp_23_16), .i_b(w_pp_24_15), .i_c(w_pp_25_14), .ow_sum(w_sum_39_39), .ow_carry(w_carry_39_39));
wire w_sum_39_37, w_carry_39_37;
math_adder_full FA_39_37(.i_a(w_pp_26_13), .i_b(w_pp_27_12), .i_c(w_pp_28_11), .ow_sum(w_sum_39_37), .ow_carry(w_carry_39_37));
wire w_sum_39_35, w_carry_39_35;
math_adder_full FA_39_35(.i_a(w_pp_29_10), .i_b(w_pp_30_09), .i_c(w_pp_31_08), .ow_sum(w_sum_39_35), .ow_carry(w_carry_39_35));
wire w_sum_39_33, w_carry_39_33;
math_adder_full FA_39_33(.i_a(w_carry_38_51), .i_b(w_carry_38_49), .i_c(w_carry_38_47), .ow_sum(w_sum_39_33), .ow_carry(w_carry_39_33));
wire w_sum_39_31, w_carry_39_31;
math_adder_full FA_39_31(.i_a(w_carry_38_45), .i_b(w_carry_38_43), .i_c(w_carry_38_41), .ow_sum(w_sum_39_31), .ow_carry(w_carry_39_31));
wire w_sum_39_29, w_carry_39_29;
math_adder_full FA_39_29(.i_a(w_carry_38_39), .i_b(w_carry_38_37), .i_c(w_carry_38_35), .ow_sum(w_sum_39_29), .ow_carry(w_carry_39_29));
wire w_sum_39_27, w_carry_39_27;
math_adder_full FA_39_27(.i_a(w_carry_38_33), .i_b(w_carry_38_31), .i_c(w_carry_38_29), .ow_sum(w_sum_39_27), .ow_carry(w_carry_39_27));
wire w_sum_39_25, w_carry_39_25;
math_adder_full FA_39_25(.i_a(w_carry_38_27), .i_b(w_carry_38_25), .i_c(w_carry_38_23), .ow_sum(w_sum_39_25), .ow_carry(w_carry_39_25));
wire w_sum_39_23, w_carry_39_23;
math_adder_full FA_39_23(.i_a(w_carry_38_21), .i_b(w_carry_38_19), .i_c(w_carry_38_17), .ow_sum(w_sum_39_23), .ow_carry(w_carry_39_23));
wire w_sum_39_21, w_carry_39_21;
math_adder_full FA_39_21(.i_a(w_carry_38_15), .i_b(w_carry_38_13), .i_c(w_carry_38_11), .ow_sum(w_sum_39_21), .ow_carry(w_carry_39_21));
wire w_sum_39_19, w_carry_39_19;
math_adder_full FA_39_19(.i_a(w_carry_38_09), .i_b(w_carry_38_07), .i_c(w_carry_38_05), .ow_sum(w_sum_39_19), .ow_carry(w_carry_39_19));
wire w_sum_39_17, w_carry_39_17;
math_adder_full FA_39_17(.i_a(w_carry_38_03), .i_b(w_sum_39_49), .i_c(w_sum_39_47), .ow_sum(w_sum_39_17), .ow_carry(w_carry_39_17));
wire w_sum_39_15, w_carry_39_15;
math_adder_full FA_39_15(.i_a(w_sum_39_45), .i_b(w_sum_39_43), .i_c(w_sum_39_41), .ow_sum(w_sum_39_15), .ow_carry(w_carry_39_15));
wire w_sum_39_13, w_carry_39_13;
math_adder_full FA_39_13(.i_a(w_sum_39_39), .i_b(w_sum_39_37), .i_c(w_sum_39_35), .ow_sum(w_sum_39_13), .ow_carry(w_carry_39_13));
wire w_sum_39_11, w_carry_39_11;
math_adder_full FA_39_11(.i_a(w_sum_39_33), .i_b(w_sum_39_31), .i_c(w_sum_39_29), .ow_sum(w_sum_39_11), .ow_carry(w_carry_39_11));
wire w_sum_39_09, w_carry_39_09;
math_adder_full FA_39_09(.i_a(w_sum_39_27), .i_b(w_sum_39_25), .i_c(w_sum_39_23), .ow_sum(w_sum_39_09), .ow_carry(w_carry_39_09));
wire w_sum_39_07, w_carry_39_07;
math_adder_full FA_39_07(.i_a(w_sum_39_21), .i_b(w_sum_39_19), .i_c(w_sum_39_17), .ow_sum(w_sum_39_07), .ow_carry(w_carry_39_07));
wire w_sum_39_05, w_carry_39_05;
math_adder_full FA_39_05(.i_a(w_sum_39_15), .i_b(w_sum_39_13), .i_c(w_sum_39_11), .ow_sum(w_sum_39_05), .ow_carry(w_carry_39_05));
wire w_sum_39_03, w_carry_39_03;
math_adder_full FA_39_03(.i_a(w_sum_39_09), .i_b(w_sum_39_07), .i_c(w_sum_39_05), .ow_sum(w_sum_39_03), .ow_carry(w_carry_39_03));
wire w_sum_40_47, w_carry_40_47;
math_adder_full FA_40_47(.i_a(w_pp_09_31), .i_b(w_pp_10_30), .i_c(w_pp_11_29), .ow_sum(w_sum_40_47), .ow_carry(w_carry_40_47));
wire w_sum_40_45, w_carry_40_45;
math_adder_full FA_40_45(.i_a(w_pp_12_28), .i_b(w_pp_13_27), .i_c(w_pp_14_26), .ow_sum(w_sum_40_45), .ow_carry(w_carry_40_45));
wire w_sum_40_43, w_carry_40_43;
math_adder_full FA_40_43(.i_a(w_pp_15_25), .i_b(w_pp_16_24), .i_c(w_pp_17_23), .ow_sum(w_sum_40_43), .ow_carry(w_carry_40_43));
wire w_sum_40_41, w_carry_40_41;
math_adder_full FA_40_41(.i_a(w_pp_18_22), .i_b(w_pp_19_21), .i_c(w_pp_20_20), .ow_sum(w_sum_40_41), .ow_carry(w_carry_40_41));
wire w_sum_40_39, w_carry_40_39;
math_adder_full FA_40_39(.i_a(w_pp_21_19), .i_b(w_pp_22_18), .i_c(w_pp_23_17), .ow_sum(w_sum_40_39), .ow_carry(w_carry_40_39));
wire w_sum_40_37, w_carry_40_37;
math_adder_full FA_40_37(.i_a(w_pp_24_16), .i_b(w_pp_25_15), .i_c(w_pp_26_14), .ow_sum(w_sum_40_37), .ow_carry(w_carry_40_37));
wire w_sum_40_35, w_carry_40_35;
math_adder_full FA_40_35(.i_a(w_pp_27_13), .i_b(w_pp_28_12), .i_c(w_pp_29_11), .ow_sum(w_sum_40_35), .ow_carry(w_carry_40_35));
wire w_sum_40_33, w_carry_40_33;
math_adder_full FA_40_33(.i_a(w_pp_30_10), .i_b(w_pp_31_09), .i_c(w_carry_39_49), .ow_sum(w_sum_40_33), .ow_carry(w_carry_40_33));
wire w_sum_40_31, w_carry_40_31;
math_adder_full FA_40_31(.i_a(w_carry_39_47), .i_b(w_carry_39_45), .i_c(w_carry_39_43), .ow_sum(w_sum_40_31), .ow_carry(w_carry_40_31));
wire w_sum_40_29, w_carry_40_29;
math_adder_full FA_40_29(.i_a(w_carry_39_41), .i_b(w_carry_39_39), .i_c(w_carry_39_37), .ow_sum(w_sum_40_29), .ow_carry(w_carry_40_29));
wire w_sum_40_27, w_carry_40_27;
math_adder_full FA_40_27(.i_a(w_carry_39_35), .i_b(w_carry_39_33), .i_c(w_carry_39_31), .ow_sum(w_sum_40_27), .ow_carry(w_carry_40_27));
wire w_sum_40_25, w_carry_40_25;
math_adder_full FA_40_25(.i_a(w_carry_39_29), .i_b(w_carry_39_27), .i_c(w_carry_39_25), .ow_sum(w_sum_40_25), .ow_carry(w_carry_40_25));
wire w_sum_40_23, w_carry_40_23;
math_adder_full FA_40_23(.i_a(w_carry_39_23), .i_b(w_carry_39_21), .i_c(w_carry_39_19), .ow_sum(w_sum_40_23), .ow_carry(w_carry_40_23));
wire w_sum_40_21, w_carry_40_21;
math_adder_full FA_40_21(.i_a(w_carry_39_17), .i_b(w_carry_39_15), .i_c(w_carry_39_13), .ow_sum(w_sum_40_21), .ow_carry(w_carry_40_21));
wire w_sum_40_19, w_carry_40_19;
math_adder_full FA_40_19(.i_a(w_carry_39_11), .i_b(w_carry_39_09), .i_c(w_carry_39_07), .ow_sum(w_sum_40_19), .ow_carry(w_carry_40_19));
wire w_sum_40_17, w_carry_40_17;
math_adder_full FA_40_17(.i_a(w_carry_39_05), .i_b(w_carry_39_03), .i_c(w_sum_40_47), .ow_sum(w_sum_40_17), .ow_carry(w_carry_40_17));
wire w_sum_40_15, w_carry_40_15;
math_adder_full FA_40_15(.i_a(w_sum_40_45), .i_b(w_sum_40_43), .i_c(w_sum_40_41), .ow_sum(w_sum_40_15), .ow_carry(w_carry_40_15));
wire w_sum_40_13, w_carry_40_13;
math_adder_full FA_40_13(.i_a(w_sum_40_39), .i_b(w_sum_40_37), .i_c(w_sum_40_35), .ow_sum(w_sum_40_13), .ow_carry(w_carry_40_13));
wire w_sum_40_11, w_carry_40_11;
math_adder_full FA_40_11(.i_a(w_sum_40_33), .i_b(w_sum_40_31), .i_c(w_sum_40_29), .ow_sum(w_sum_40_11), .ow_carry(w_carry_40_11));
wire w_sum_40_09, w_carry_40_09;
math_adder_full FA_40_09(.i_a(w_sum_40_27), .i_b(w_sum_40_25), .i_c(w_sum_40_23), .ow_sum(w_sum_40_09), .ow_carry(w_carry_40_09));
wire w_sum_40_07, w_carry_40_07;
math_adder_full FA_40_07(.i_a(w_sum_40_21), .i_b(w_sum_40_19), .i_c(w_sum_40_17), .ow_sum(w_sum_40_07), .ow_carry(w_carry_40_07));
wire w_sum_40_05, w_carry_40_05;
math_adder_full FA_40_05(.i_a(w_sum_40_15), .i_b(w_sum_40_13), .i_c(w_sum_40_11), .ow_sum(w_sum_40_05), .ow_carry(w_carry_40_05));
wire w_sum_40_03, w_carry_40_03;
math_adder_full FA_40_03(.i_a(w_sum_40_09), .i_b(w_sum_40_07), .i_c(w_sum_40_05), .ow_sum(w_sum_40_03), .ow_carry(w_carry_40_03));
wire w_sum_41_45, w_carry_41_45;
math_adder_full FA_41_45(.i_a(w_pp_10_31), .i_b(w_pp_11_30), .i_c(w_pp_12_29), .ow_sum(w_sum_41_45), .ow_carry(w_carry_41_45));
wire w_sum_41_43, w_carry_41_43;
math_adder_full FA_41_43(.i_a(w_pp_13_28), .i_b(w_pp_14_27), .i_c(w_pp_15_26), .ow_sum(w_sum_41_43), .ow_carry(w_carry_41_43));
wire w_sum_41_41, w_carry_41_41;
math_adder_full FA_41_41(.i_a(w_pp_16_25), .i_b(w_pp_17_24), .i_c(w_pp_18_23), .ow_sum(w_sum_41_41), .ow_carry(w_carry_41_41));
wire w_sum_41_39, w_carry_41_39;
math_adder_full FA_41_39(.i_a(w_pp_19_22), .i_b(w_pp_20_21), .i_c(w_pp_21_20), .ow_sum(w_sum_41_39), .ow_carry(w_carry_41_39));
wire w_sum_41_37, w_carry_41_37;
math_adder_full FA_41_37(.i_a(w_pp_22_19), .i_b(w_pp_23_18), .i_c(w_pp_24_17), .ow_sum(w_sum_41_37), .ow_carry(w_carry_41_37));
wire w_sum_41_35, w_carry_41_35;
math_adder_full FA_41_35(.i_a(w_pp_25_16), .i_b(w_pp_26_15), .i_c(w_pp_27_14), .ow_sum(w_sum_41_35), .ow_carry(w_carry_41_35));
wire w_sum_41_33, w_carry_41_33;
math_adder_full FA_41_33(.i_a(w_pp_28_13), .i_b(w_pp_29_12), .i_c(w_pp_30_11), .ow_sum(w_sum_41_33), .ow_carry(w_carry_41_33));
wire w_sum_41_31, w_carry_41_31;
math_adder_full FA_41_31(.i_a(w_pp_31_10), .i_b(w_carry_40_47), .i_c(w_carry_40_45), .ow_sum(w_sum_41_31), .ow_carry(w_carry_41_31));
wire w_sum_41_29, w_carry_41_29;
math_adder_full FA_41_29(.i_a(w_carry_40_43), .i_b(w_carry_40_41), .i_c(w_carry_40_39), .ow_sum(w_sum_41_29), .ow_carry(w_carry_41_29));
wire w_sum_41_27, w_carry_41_27;
math_adder_full FA_41_27(.i_a(w_carry_40_37), .i_b(w_carry_40_35), .i_c(w_carry_40_33), .ow_sum(w_sum_41_27), .ow_carry(w_carry_41_27));
wire w_sum_41_25, w_carry_41_25;
math_adder_full FA_41_25(.i_a(w_carry_40_31), .i_b(w_carry_40_29), .i_c(w_carry_40_27), .ow_sum(w_sum_41_25), .ow_carry(w_carry_41_25));
wire w_sum_41_23, w_carry_41_23;
math_adder_full FA_41_23(.i_a(w_carry_40_25), .i_b(w_carry_40_23), .i_c(w_carry_40_21), .ow_sum(w_sum_41_23), .ow_carry(w_carry_41_23));
wire w_sum_41_21, w_carry_41_21;
math_adder_full FA_41_21(.i_a(w_carry_40_19), .i_b(w_carry_40_17), .i_c(w_carry_40_15), .ow_sum(w_sum_41_21), .ow_carry(w_carry_41_21));
wire w_sum_41_19, w_carry_41_19;
math_adder_full FA_41_19(.i_a(w_carry_40_13), .i_b(w_carry_40_11), .i_c(w_carry_40_09), .ow_sum(w_sum_41_19), .ow_carry(w_carry_41_19));
wire w_sum_41_17, w_carry_41_17;
math_adder_full FA_41_17(.i_a(w_carry_40_07), .i_b(w_carry_40_05), .i_c(w_carry_40_03), .ow_sum(w_sum_41_17), .ow_carry(w_carry_41_17));
wire w_sum_41_15, w_carry_41_15;
math_adder_full FA_41_15(.i_a(w_sum_41_45), .i_b(w_sum_41_43), .i_c(w_sum_41_41), .ow_sum(w_sum_41_15), .ow_carry(w_carry_41_15));
wire w_sum_41_13, w_carry_41_13;
math_adder_full FA_41_13(.i_a(w_sum_41_39), .i_b(w_sum_41_37), .i_c(w_sum_41_35), .ow_sum(w_sum_41_13), .ow_carry(w_carry_41_13));
wire w_sum_41_11, w_carry_41_11;
math_adder_full FA_41_11(.i_a(w_sum_41_33), .i_b(w_sum_41_31), .i_c(w_sum_41_29), .ow_sum(w_sum_41_11), .ow_carry(w_carry_41_11));
wire w_sum_41_09, w_carry_41_09;
math_adder_full FA_41_09(.i_a(w_sum_41_27), .i_b(w_sum_41_25), .i_c(w_sum_41_23), .ow_sum(w_sum_41_09), .ow_carry(w_carry_41_09));
wire w_sum_41_07, w_carry_41_07;
math_adder_full FA_41_07(.i_a(w_sum_41_21), .i_b(w_sum_41_19), .i_c(w_sum_41_17), .ow_sum(w_sum_41_07), .ow_carry(w_carry_41_07));
wire w_sum_41_05, w_carry_41_05;
math_adder_full FA_41_05(.i_a(w_sum_41_15), .i_b(w_sum_41_13), .i_c(w_sum_41_11), .ow_sum(w_sum_41_05), .ow_carry(w_carry_41_05));
wire w_sum_41_03, w_carry_41_03;
math_adder_full FA_41_03(.i_a(w_sum_41_09), .i_b(w_sum_41_07), .i_c(w_sum_41_05), .ow_sum(w_sum_41_03), .ow_carry(w_carry_41_03));
wire w_sum_42_43, w_carry_42_43;
math_adder_full FA_42_43(.i_a(w_pp_11_31), .i_b(w_pp_12_30), .i_c(w_pp_13_29), .ow_sum(w_sum_42_43), .ow_carry(w_carry_42_43));
wire w_sum_42_41, w_carry_42_41;
math_adder_full FA_42_41(.i_a(w_pp_14_28), .i_b(w_pp_15_27), .i_c(w_pp_16_26), .ow_sum(w_sum_42_41), .ow_carry(w_carry_42_41));
wire w_sum_42_39, w_carry_42_39;
math_adder_full FA_42_39(.i_a(w_pp_17_25), .i_b(w_pp_18_24), .i_c(w_pp_19_23), .ow_sum(w_sum_42_39), .ow_carry(w_carry_42_39));
wire w_sum_42_37, w_carry_42_37;
math_adder_full FA_42_37(.i_a(w_pp_20_22), .i_b(w_pp_21_21), .i_c(w_pp_22_20), .ow_sum(w_sum_42_37), .ow_carry(w_carry_42_37));
wire w_sum_42_35, w_carry_42_35;
math_adder_full FA_42_35(.i_a(w_pp_23_19), .i_b(w_pp_24_18), .i_c(w_pp_25_17), .ow_sum(w_sum_42_35), .ow_carry(w_carry_42_35));
wire w_sum_42_33, w_carry_42_33;
math_adder_full FA_42_33(.i_a(w_pp_26_16), .i_b(w_pp_27_15), .i_c(w_pp_28_14), .ow_sum(w_sum_42_33), .ow_carry(w_carry_42_33));
wire w_sum_42_31, w_carry_42_31;
math_adder_full FA_42_31(.i_a(w_pp_29_13), .i_b(w_pp_30_12), .i_c(w_pp_31_11), .ow_sum(w_sum_42_31), .ow_carry(w_carry_42_31));
wire w_sum_42_29, w_carry_42_29;
math_adder_full FA_42_29(.i_a(w_carry_41_45), .i_b(w_carry_41_43), .i_c(w_carry_41_41), .ow_sum(w_sum_42_29), .ow_carry(w_carry_42_29));
wire w_sum_42_27, w_carry_42_27;
math_adder_full FA_42_27(.i_a(w_carry_41_39), .i_b(w_carry_41_37), .i_c(w_carry_41_35), .ow_sum(w_sum_42_27), .ow_carry(w_carry_42_27));
wire w_sum_42_25, w_carry_42_25;
math_adder_full FA_42_25(.i_a(w_carry_41_33), .i_b(w_carry_41_31), .i_c(w_carry_41_29), .ow_sum(w_sum_42_25), .ow_carry(w_carry_42_25));
wire w_sum_42_23, w_carry_42_23;
math_adder_full FA_42_23(.i_a(w_carry_41_27), .i_b(w_carry_41_25), .i_c(w_carry_41_23), .ow_sum(w_sum_42_23), .ow_carry(w_carry_42_23));
wire w_sum_42_21, w_carry_42_21;
math_adder_full FA_42_21(.i_a(w_carry_41_21), .i_b(w_carry_41_19), .i_c(w_carry_41_17), .ow_sum(w_sum_42_21), .ow_carry(w_carry_42_21));
wire w_sum_42_19, w_carry_42_19;
math_adder_full FA_42_19(.i_a(w_carry_41_15), .i_b(w_carry_41_13), .i_c(w_carry_41_11), .ow_sum(w_sum_42_19), .ow_carry(w_carry_42_19));
wire w_sum_42_17, w_carry_42_17;
math_adder_full FA_42_17(.i_a(w_carry_41_09), .i_b(w_carry_41_07), .i_c(w_carry_41_05), .ow_sum(w_sum_42_17), .ow_carry(w_carry_42_17));
wire w_sum_42_15, w_carry_42_15;
math_adder_full FA_42_15(.i_a(w_carry_41_03), .i_b(w_sum_42_43), .i_c(w_sum_42_41), .ow_sum(w_sum_42_15), .ow_carry(w_carry_42_15));
wire w_sum_42_13, w_carry_42_13;
math_adder_full FA_42_13(.i_a(w_sum_42_39), .i_b(w_sum_42_37), .i_c(w_sum_42_35), .ow_sum(w_sum_42_13), .ow_carry(w_carry_42_13));
wire w_sum_42_11, w_carry_42_11;
math_adder_full FA_42_11(.i_a(w_sum_42_33), .i_b(w_sum_42_31), .i_c(w_sum_42_29), .ow_sum(w_sum_42_11), .ow_carry(w_carry_42_11));
wire w_sum_42_09, w_carry_42_09;
math_adder_full FA_42_09(.i_a(w_sum_42_27), .i_b(w_sum_42_25), .i_c(w_sum_42_23), .ow_sum(w_sum_42_09), .ow_carry(w_carry_42_09));
wire w_sum_42_07, w_carry_42_07;
math_adder_full FA_42_07(.i_a(w_sum_42_21), .i_b(w_sum_42_19), .i_c(w_sum_42_17), .ow_sum(w_sum_42_07), .ow_carry(w_carry_42_07));
wire w_sum_42_05, w_carry_42_05;
math_adder_full FA_42_05(.i_a(w_sum_42_15), .i_b(w_sum_42_13), .i_c(w_sum_42_11), .ow_sum(w_sum_42_05), .ow_carry(w_carry_42_05));
wire w_sum_42_03, w_carry_42_03;
math_adder_full FA_42_03(.i_a(w_sum_42_09), .i_b(w_sum_42_07), .i_c(w_sum_42_05), .ow_sum(w_sum_42_03), .ow_carry(w_carry_42_03));
wire w_sum_43_41, w_carry_43_41;
math_adder_full FA_43_41(.i_a(w_pp_12_31), .i_b(w_pp_13_30), .i_c(w_pp_14_29), .ow_sum(w_sum_43_41), .ow_carry(w_carry_43_41));
wire w_sum_43_39, w_carry_43_39;
math_adder_full FA_43_39(.i_a(w_pp_15_28), .i_b(w_pp_16_27), .i_c(w_pp_17_26), .ow_sum(w_sum_43_39), .ow_carry(w_carry_43_39));
wire w_sum_43_37, w_carry_43_37;
math_adder_full FA_43_37(.i_a(w_pp_18_25), .i_b(w_pp_19_24), .i_c(w_pp_20_23), .ow_sum(w_sum_43_37), .ow_carry(w_carry_43_37));
wire w_sum_43_35, w_carry_43_35;
math_adder_full FA_43_35(.i_a(w_pp_21_22), .i_b(w_pp_22_21), .i_c(w_pp_23_20), .ow_sum(w_sum_43_35), .ow_carry(w_carry_43_35));
wire w_sum_43_33, w_carry_43_33;
math_adder_full FA_43_33(.i_a(w_pp_24_19), .i_b(w_pp_25_18), .i_c(w_pp_26_17), .ow_sum(w_sum_43_33), .ow_carry(w_carry_43_33));
wire w_sum_43_31, w_carry_43_31;
math_adder_full FA_43_31(.i_a(w_pp_27_16), .i_b(w_pp_28_15), .i_c(w_pp_29_14), .ow_sum(w_sum_43_31), .ow_carry(w_carry_43_31));
wire w_sum_43_29, w_carry_43_29;
math_adder_full FA_43_29(.i_a(w_pp_30_13), .i_b(w_pp_31_12), .i_c(w_carry_42_43), .ow_sum(w_sum_43_29), .ow_carry(w_carry_43_29));
wire w_sum_43_27, w_carry_43_27;
math_adder_full FA_43_27(.i_a(w_carry_42_41), .i_b(w_carry_42_39), .i_c(w_carry_42_37), .ow_sum(w_sum_43_27), .ow_carry(w_carry_43_27));
wire w_sum_43_25, w_carry_43_25;
math_adder_full FA_43_25(.i_a(w_carry_42_35), .i_b(w_carry_42_33), .i_c(w_carry_42_31), .ow_sum(w_sum_43_25), .ow_carry(w_carry_43_25));
wire w_sum_43_23, w_carry_43_23;
math_adder_full FA_43_23(.i_a(w_carry_42_29), .i_b(w_carry_42_27), .i_c(w_carry_42_25), .ow_sum(w_sum_43_23), .ow_carry(w_carry_43_23));
wire w_sum_43_21, w_carry_43_21;
math_adder_full FA_43_21(.i_a(w_carry_42_23), .i_b(w_carry_42_21), .i_c(w_carry_42_19), .ow_sum(w_sum_43_21), .ow_carry(w_carry_43_21));
wire w_sum_43_19, w_carry_43_19;
math_adder_full FA_43_19(.i_a(w_carry_42_17), .i_b(w_carry_42_15), .i_c(w_carry_42_13), .ow_sum(w_sum_43_19), .ow_carry(w_carry_43_19));
wire w_sum_43_17, w_carry_43_17;
math_adder_full FA_43_17(.i_a(w_carry_42_11), .i_b(w_carry_42_09), .i_c(w_carry_42_07), .ow_sum(w_sum_43_17), .ow_carry(w_carry_43_17));
wire w_sum_43_15, w_carry_43_15;
math_adder_full FA_43_15(.i_a(w_carry_42_05), .i_b(w_carry_42_03), .i_c(w_sum_43_41), .ow_sum(w_sum_43_15), .ow_carry(w_carry_43_15));
wire w_sum_43_13, w_carry_43_13;
math_adder_full FA_43_13(.i_a(w_sum_43_39), .i_b(w_sum_43_37), .i_c(w_sum_43_35), .ow_sum(w_sum_43_13), .ow_carry(w_carry_43_13));
wire w_sum_43_11, w_carry_43_11;
math_adder_full FA_43_11(.i_a(w_sum_43_33), .i_b(w_sum_43_31), .i_c(w_sum_43_29), .ow_sum(w_sum_43_11), .ow_carry(w_carry_43_11));
wire w_sum_43_09, w_carry_43_09;
math_adder_full FA_43_09(.i_a(w_sum_43_27), .i_b(w_sum_43_25), .i_c(w_sum_43_23), .ow_sum(w_sum_43_09), .ow_carry(w_carry_43_09));
wire w_sum_43_07, w_carry_43_07;
math_adder_full FA_43_07(.i_a(w_sum_43_21), .i_b(w_sum_43_19), .i_c(w_sum_43_17), .ow_sum(w_sum_43_07), .ow_carry(w_carry_43_07));
wire w_sum_43_05, w_carry_43_05;
math_adder_full FA_43_05(.i_a(w_sum_43_15), .i_b(w_sum_43_13), .i_c(w_sum_43_11), .ow_sum(w_sum_43_05), .ow_carry(w_carry_43_05));
wire w_sum_43_03, w_carry_43_03;
math_adder_full FA_43_03(.i_a(w_sum_43_09), .i_b(w_sum_43_07), .i_c(w_sum_43_05), .ow_sum(w_sum_43_03), .ow_carry(w_carry_43_03));
wire w_sum_44_39, w_carry_44_39;
math_adder_full FA_44_39(.i_a(w_pp_13_31), .i_b(w_pp_14_30), .i_c(w_pp_15_29), .ow_sum(w_sum_44_39), .ow_carry(w_carry_44_39));
wire w_sum_44_37, w_carry_44_37;
math_adder_full FA_44_37(.i_a(w_pp_16_28), .i_b(w_pp_17_27), .i_c(w_pp_18_26), .ow_sum(w_sum_44_37), .ow_carry(w_carry_44_37));
wire w_sum_44_35, w_carry_44_35;
math_adder_full FA_44_35(.i_a(w_pp_19_25), .i_b(w_pp_20_24), .i_c(w_pp_21_23), .ow_sum(w_sum_44_35), .ow_carry(w_carry_44_35));
wire w_sum_44_33, w_carry_44_33;
math_adder_full FA_44_33(.i_a(w_pp_22_22), .i_b(w_pp_23_21), .i_c(w_pp_24_20), .ow_sum(w_sum_44_33), .ow_carry(w_carry_44_33));
wire w_sum_44_31, w_carry_44_31;
math_adder_full FA_44_31(.i_a(w_pp_25_19), .i_b(w_pp_26_18), .i_c(w_pp_27_17), .ow_sum(w_sum_44_31), .ow_carry(w_carry_44_31));
wire w_sum_44_29, w_carry_44_29;
math_adder_full FA_44_29(.i_a(w_pp_28_16), .i_b(w_pp_29_15), .i_c(w_pp_30_14), .ow_sum(w_sum_44_29), .ow_carry(w_carry_44_29));
wire w_sum_44_27, w_carry_44_27;
math_adder_full FA_44_27(.i_a(w_pp_31_13), .i_b(w_carry_43_41), .i_c(w_carry_43_39), .ow_sum(w_sum_44_27), .ow_carry(w_carry_44_27));
wire w_sum_44_25, w_carry_44_25;
math_adder_full FA_44_25(.i_a(w_carry_43_37), .i_b(w_carry_43_35), .i_c(w_carry_43_33), .ow_sum(w_sum_44_25), .ow_carry(w_carry_44_25));
wire w_sum_44_23, w_carry_44_23;
math_adder_full FA_44_23(.i_a(w_carry_43_31), .i_b(w_carry_43_29), .i_c(w_carry_43_27), .ow_sum(w_sum_44_23), .ow_carry(w_carry_44_23));
wire w_sum_44_21, w_carry_44_21;
math_adder_full FA_44_21(.i_a(w_carry_43_25), .i_b(w_carry_43_23), .i_c(w_carry_43_21), .ow_sum(w_sum_44_21), .ow_carry(w_carry_44_21));
wire w_sum_44_19, w_carry_44_19;
math_adder_full FA_44_19(.i_a(w_carry_43_19), .i_b(w_carry_43_17), .i_c(w_carry_43_15), .ow_sum(w_sum_44_19), .ow_carry(w_carry_44_19));
wire w_sum_44_17, w_carry_44_17;
math_adder_full FA_44_17(.i_a(w_carry_43_13), .i_b(w_carry_43_11), .i_c(w_carry_43_09), .ow_sum(w_sum_44_17), .ow_carry(w_carry_44_17));
wire w_sum_44_15, w_carry_44_15;
math_adder_full FA_44_15(.i_a(w_carry_43_07), .i_b(w_carry_43_05), .i_c(w_carry_43_03), .ow_sum(w_sum_44_15), .ow_carry(w_carry_44_15));
wire w_sum_44_13, w_carry_44_13;
math_adder_full FA_44_13(.i_a(w_sum_44_39), .i_b(w_sum_44_37), .i_c(w_sum_44_35), .ow_sum(w_sum_44_13), .ow_carry(w_carry_44_13));
wire w_sum_44_11, w_carry_44_11;
math_adder_full FA_44_11(.i_a(w_sum_44_33), .i_b(w_sum_44_31), .i_c(w_sum_44_29), .ow_sum(w_sum_44_11), .ow_carry(w_carry_44_11));
wire w_sum_44_09, w_carry_44_09;
math_adder_full FA_44_09(.i_a(w_sum_44_27), .i_b(w_sum_44_25), .i_c(w_sum_44_23), .ow_sum(w_sum_44_09), .ow_carry(w_carry_44_09));
wire w_sum_44_07, w_carry_44_07;
math_adder_full FA_44_07(.i_a(w_sum_44_21), .i_b(w_sum_44_19), .i_c(w_sum_44_17), .ow_sum(w_sum_44_07), .ow_carry(w_carry_44_07));
wire w_sum_44_05, w_carry_44_05;
math_adder_full FA_44_05(.i_a(w_sum_44_15), .i_b(w_sum_44_13), .i_c(w_sum_44_11), .ow_sum(w_sum_44_05), .ow_carry(w_carry_44_05));
wire w_sum_44_03, w_carry_44_03;
math_adder_full FA_44_03(.i_a(w_sum_44_09), .i_b(w_sum_44_07), .i_c(w_sum_44_05), .ow_sum(w_sum_44_03), .ow_carry(w_carry_44_03));
wire w_sum_45_37, w_carry_45_37;
math_adder_full FA_45_37(.i_a(w_pp_14_31), .i_b(w_pp_15_30), .i_c(w_pp_16_29), .ow_sum(w_sum_45_37), .ow_carry(w_carry_45_37));
wire w_sum_45_35, w_carry_45_35;
math_adder_full FA_45_35(.i_a(w_pp_17_28), .i_b(w_pp_18_27), .i_c(w_pp_19_26), .ow_sum(w_sum_45_35), .ow_carry(w_carry_45_35));
wire w_sum_45_33, w_carry_45_33;
math_adder_full FA_45_33(.i_a(w_pp_20_25), .i_b(w_pp_21_24), .i_c(w_pp_22_23), .ow_sum(w_sum_45_33), .ow_carry(w_carry_45_33));
wire w_sum_45_31, w_carry_45_31;
math_adder_full FA_45_31(.i_a(w_pp_23_22), .i_b(w_pp_24_21), .i_c(w_pp_25_20), .ow_sum(w_sum_45_31), .ow_carry(w_carry_45_31));
wire w_sum_45_29, w_carry_45_29;
math_adder_full FA_45_29(.i_a(w_pp_26_19), .i_b(w_pp_27_18), .i_c(w_pp_28_17), .ow_sum(w_sum_45_29), .ow_carry(w_carry_45_29));
wire w_sum_45_27, w_carry_45_27;
math_adder_full FA_45_27(.i_a(w_pp_29_16), .i_b(w_pp_30_15), .i_c(w_pp_31_14), .ow_sum(w_sum_45_27), .ow_carry(w_carry_45_27));
wire w_sum_45_25, w_carry_45_25;
math_adder_full FA_45_25(.i_a(w_carry_44_39), .i_b(w_carry_44_37), .i_c(w_carry_44_35), .ow_sum(w_sum_45_25), .ow_carry(w_carry_45_25));
wire w_sum_45_23, w_carry_45_23;
math_adder_full FA_45_23(.i_a(w_carry_44_33), .i_b(w_carry_44_31), .i_c(w_carry_44_29), .ow_sum(w_sum_45_23), .ow_carry(w_carry_45_23));
wire w_sum_45_21, w_carry_45_21;
math_adder_full FA_45_21(.i_a(w_carry_44_27), .i_b(w_carry_44_25), .i_c(w_carry_44_23), .ow_sum(w_sum_45_21), .ow_carry(w_carry_45_21));
wire w_sum_45_19, w_carry_45_19;
math_adder_full FA_45_19(.i_a(w_carry_44_21), .i_b(w_carry_44_19), .i_c(w_carry_44_17), .ow_sum(w_sum_45_19), .ow_carry(w_carry_45_19));
wire w_sum_45_17, w_carry_45_17;
math_adder_full FA_45_17(.i_a(w_carry_44_15), .i_b(w_carry_44_13), .i_c(w_carry_44_11), .ow_sum(w_sum_45_17), .ow_carry(w_carry_45_17));
wire w_sum_45_15, w_carry_45_15;
math_adder_full FA_45_15(.i_a(w_carry_44_09), .i_b(w_carry_44_07), .i_c(w_carry_44_05), .ow_sum(w_sum_45_15), .ow_carry(w_carry_45_15));
wire w_sum_45_13, w_carry_45_13;
math_adder_full FA_45_13(.i_a(w_carry_44_03), .i_b(w_sum_45_37), .i_c(w_sum_45_35), .ow_sum(w_sum_45_13), .ow_carry(w_carry_45_13));
wire w_sum_45_11, w_carry_45_11;
math_adder_full FA_45_11(.i_a(w_sum_45_33), .i_b(w_sum_45_31), .i_c(w_sum_45_29), .ow_sum(w_sum_45_11), .ow_carry(w_carry_45_11));
wire w_sum_45_09, w_carry_45_09;
math_adder_full FA_45_09(.i_a(w_sum_45_27), .i_b(w_sum_45_25), .i_c(w_sum_45_23), .ow_sum(w_sum_45_09), .ow_carry(w_carry_45_09));
wire w_sum_45_07, w_carry_45_07;
math_adder_full FA_45_07(.i_a(w_sum_45_21), .i_b(w_sum_45_19), .i_c(w_sum_45_17), .ow_sum(w_sum_45_07), .ow_carry(w_carry_45_07));
wire w_sum_45_05, w_carry_45_05;
math_adder_full FA_45_05(.i_a(w_sum_45_15), .i_b(w_sum_45_13), .i_c(w_sum_45_11), .ow_sum(w_sum_45_05), .ow_carry(w_carry_45_05));
wire w_sum_45_03, w_carry_45_03;
math_adder_full FA_45_03(.i_a(w_sum_45_09), .i_b(w_sum_45_07), .i_c(w_sum_45_05), .ow_sum(w_sum_45_03), .ow_carry(w_carry_45_03));
wire w_sum_46_35, w_carry_46_35;
math_adder_full FA_46_35(.i_a(w_pp_15_31), .i_b(w_pp_16_30), .i_c(w_pp_17_29), .ow_sum(w_sum_46_35), .ow_carry(w_carry_46_35));
wire w_sum_46_33, w_carry_46_33;
math_adder_full FA_46_33(.i_a(w_pp_18_28), .i_b(w_pp_19_27), .i_c(w_pp_20_26), .ow_sum(w_sum_46_33), .ow_carry(w_carry_46_33));
wire w_sum_46_31, w_carry_46_31;
math_adder_full FA_46_31(.i_a(w_pp_21_25), .i_b(w_pp_22_24), .i_c(w_pp_23_23), .ow_sum(w_sum_46_31), .ow_carry(w_carry_46_31));
wire w_sum_46_29, w_carry_46_29;
math_adder_full FA_46_29(.i_a(w_pp_24_22), .i_b(w_pp_25_21), .i_c(w_pp_26_20), .ow_sum(w_sum_46_29), .ow_carry(w_carry_46_29));
wire w_sum_46_27, w_carry_46_27;
math_adder_full FA_46_27(.i_a(w_pp_27_19), .i_b(w_pp_28_18), .i_c(w_pp_29_17), .ow_sum(w_sum_46_27), .ow_carry(w_carry_46_27));
wire w_sum_46_25, w_carry_46_25;
math_adder_full FA_46_25(.i_a(w_pp_30_16), .i_b(w_pp_31_15), .i_c(w_carry_45_37), .ow_sum(w_sum_46_25), .ow_carry(w_carry_46_25));
wire w_sum_46_23, w_carry_46_23;
math_adder_full FA_46_23(.i_a(w_carry_45_35), .i_b(w_carry_45_33), .i_c(w_carry_45_31), .ow_sum(w_sum_46_23), .ow_carry(w_carry_46_23));
wire w_sum_46_21, w_carry_46_21;
math_adder_full FA_46_21(.i_a(w_carry_45_29), .i_b(w_carry_45_27), .i_c(w_carry_45_25), .ow_sum(w_sum_46_21), .ow_carry(w_carry_46_21));
wire w_sum_46_19, w_carry_46_19;
math_adder_full FA_46_19(.i_a(w_carry_45_23), .i_b(w_carry_45_21), .i_c(w_carry_45_19), .ow_sum(w_sum_46_19), .ow_carry(w_carry_46_19));
wire w_sum_46_17, w_carry_46_17;
math_adder_full FA_46_17(.i_a(w_carry_45_17), .i_b(w_carry_45_15), .i_c(w_carry_45_13), .ow_sum(w_sum_46_17), .ow_carry(w_carry_46_17));
wire w_sum_46_15, w_carry_46_15;
math_adder_full FA_46_15(.i_a(w_carry_45_11), .i_b(w_carry_45_09), .i_c(w_carry_45_07), .ow_sum(w_sum_46_15), .ow_carry(w_carry_46_15));
wire w_sum_46_13, w_carry_46_13;
math_adder_full FA_46_13(.i_a(w_carry_45_05), .i_b(w_carry_45_03), .i_c(w_sum_46_35), .ow_sum(w_sum_46_13), .ow_carry(w_carry_46_13));
wire w_sum_46_11, w_carry_46_11;
math_adder_full FA_46_11(.i_a(w_sum_46_33), .i_b(w_sum_46_31), .i_c(w_sum_46_29), .ow_sum(w_sum_46_11), .ow_carry(w_carry_46_11));
wire w_sum_46_09, w_carry_46_09;
math_adder_full FA_46_09(.i_a(w_sum_46_27), .i_b(w_sum_46_25), .i_c(w_sum_46_23), .ow_sum(w_sum_46_09), .ow_carry(w_carry_46_09));
wire w_sum_46_07, w_carry_46_07;
math_adder_full FA_46_07(.i_a(w_sum_46_21), .i_b(w_sum_46_19), .i_c(w_sum_46_17), .ow_sum(w_sum_46_07), .ow_carry(w_carry_46_07));
wire w_sum_46_05, w_carry_46_05;
math_adder_full FA_46_05(.i_a(w_sum_46_15), .i_b(w_sum_46_13), .i_c(w_sum_46_11), .ow_sum(w_sum_46_05), .ow_carry(w_carry_46_05));
wire w_sum_46_03, w_carry_46_03;
math_adder_full FA_46_03(.i_a(w_sum_46_09), .i_b(w_sum_46_07), .i_c(w_sum_46_05), .ow_sum(w_sum_46_03), .ow_carry(w_carry_46_03));
wire w_sum_47_33, w_carry_47_33;
math_adder_full FA_47_33(.i_a(w_pp_16_31), .i_b(w_pp_17_30), .i_c(w_pp_18_29), .ow_sum(w_sum_47_33), .ow_carry(w_carry_47_33));
wire w_sum_47_31, w_carry_47_31;
math_adder_full FA_47_31(.i_a(w_pp_19_28), .i_b(w_pp_20_27), .i_c(w_pp_21_26), .ow_sum(w_sum_47_31), .ow_carry(w_carry_47_31));
wire w_sum_47_29, w_carry_47_29;
math_adder_full FA_47_29(.i_a(w_pp_22_25), .i_b(w_pp_23_24), .i_c(w_pp_24_23), .ow_sum(w_sum_47_29), .ow_carry(w_carry_47_29));
wire w_sum_47_27, w_carry_47_27;
math_adder_full FA_47_27(.i_a(w_pp_25_22), .i_b(w_pp_26_21), .i_c(w_pp_27_20), .ow_sum(w_sum_47_27), .ow_carry(w_carry_47_27));
wire w_sum_47_25, w_carry_47_25;
math_adder_full FA_47_25(.i_a(w_pp_28_19), .i_b(w_pp_29_18), .i_c(w_pp_30_17), .ow_sum(w_sum_47_25), .ow_carry(w_carry_47_25));
wire w_sum_47_23, w_carry_47_23;
math_adder_full FA_47_23(.i_a(w_pp_31_16), .i_b(w_carry_46_35), .i_c(w_carry_46_33), .ow_sum(w_sum_47_23), .ow_carry(w_carry_47_23));
wire w_sum_47_21, w_carry_47_21;
math_adder_full FA_47_21(.i_a(w_carry_46_31), .i_b(w_carry_46_29), .i_c(w_carry_46_27), .ow_sum(w_sum_47_21), .ow_carry(w_carry_47_21));
wire w_sum_47_19, w_carry_47_19;
math_adder_full FA_47_19(.i_a(w_carry_46_25), .i_b(w_carry_46_23), .i_c(w_carry_46_21), .ow_sum(w_sum_47_19), .ow_carry(w_carry_47_19));
wire w_sum_47_17, w_carry_47_17;
math_adder_full FA_47_17(.i_a(w_carry_46_19), .i_b(w_carry_46_17), .i_c(w_carry_46_15), .ow_sum(w_sum_47_17), .ow_carry(w_carry_47_17));
wire w_sum_47_15, w_carry_47_15;
math_adder_full FA_47_15(.i_a(w_carry_46_13), .i_b(w_carry_46_11), .i_c(w_carry_46_09), .ow_sum(w_sum_47_15), .ow_carry(w_carry_47_15));
wire w_sum_47_13, w_carry_47_13;
math_adder_full FA_47_13(.i_a(w_carry_46_07), .i_b(w_carry_46_05), .i_c(w_carry_46_03), .ow_sum(w_sum_47_13), .ow_carry(w_carry_47_13));
wire w_sum_47_11, w_carry_47_11;
math_adder_full FA_47_11(.i_a(w_sum_47_33), .i_b(w_sum_47_31), .i_c(w_sum_47_29), .ow_sum(w_sum_47_11), .ow_carry(w_carry_47_11));
wire w_sum_47_09, w_carry_47_09;
math_adder_full FA_47_09(.i_a(w_sum_47_27), .i_b(w_sum_47_25), .i_c(w_sum_47_23), .ow_sum(w_sum_47_09), .ow_carry(w_carry_47_09));
wire w_sum_47_07, w_carry_47_07;
math_adder_full FA_47_07(.i_a(w_sum_47_21), .i_b(w_sum_47_19), .i_c(w_sum_47_17), .ow_sum(w_sum_47_07), .ow_carry(w_carry_47_07));
wire w_sum_47_05, w_carry_47_05;
math_adder_full FA_47_05(.i_a(w_sum_47_15), .i_b(w_sum_47_13), .i_c(w_sum_47_11), .ow_sum(w_sum_47_05), .ow_carry(w_carry_47_05));
wire w_sum_47_03, w_carry_47_03;
math_adder_full FA_47_03(.i_a(w_sum_47_09), .i_b(w_sum_47_07), .i_c(w_sum_47_05), .ow_sum(w_sum_47_03), .ow_carry(w_carry_47_03));
wire w_sum_48_31, w_carry_48_31;
math_adder_full FA_48_31(.i_a(w_pp_17_31), .i_b(w_pp_18_30), .i_c(w_pp_19_29), .ow_sum(w_sum_48_31), .ow_carry(w_carry_48_31));
wire w_sum_48_29, w_carry_48_29;
math_adder_full FA_48_29(.i_a(w_pp_20_28), .i_b(w_pp_21_27), .i_c(w_pp_22_26), .ow_sum(w_sum_48_29), .ow_carry(w_carry_48_29));
wire w_sum_48_27, w_carry_48_27;
math_adder_full FA_48_27(.i_a(w_pp_23_25), .i_b(w_pp_24_24), .i_c(w_pp_25_23), .ow_sum(w_sum_48_27), .ow_carry(w_carry_48_27));
wire w_sum_48_25, w_carry_48_25;
math_adder_full FA_48_25(.i_a(w_pp_26_22), .i_b(w_pp_27_21), .i_c(w_pp_28_20), .ow_sum(w_sum_48_25), .ow_carry(w_carry_48_25));
wire w_sum_48_23, w_carry_48_23;
math_adder_full FA_48_23(.i_a(w_pp_29_19), .i_b(w_pp_30_18), .i_c(w_pp_31_17), .ow_sum(w_sum_48_23), .ow_carry(w_carry_48_23));
wire w_sum_48_21, w_carry_48_21;
math_adder_full FA_48_21(.i_a(w_carry_47_33), .i_b(w_carry_47_31), .i_c(w_carry_47_29), .ow_sum(w_sum_48_21), .ow_carry(w_carry_48_21));
wire w_sum_48_19, w_carry_48_19;
math_adder_full FA_48_19(.i_a(w_carry_47_27), .i_b(w_carry_47_25), .i_c(w_carry_47_23), .ow_sum(w_sum_48_19), .ow_carry(w_carry_48_19));
wire w_sum_48_17, w_carry_48_17;
math_adder_full FA_48_17(.i_a(w_carry_47_21), .i_b(w_carry_47_19), .i_c(w_carry_47_17), .ow_sum(w_sum_48_17), .ow_carry(w_carry_48_17));
wire w_sum_48_15, w_carry_48_15;
math_adder_full FA_48_15(.i_a(w_carry_47_15), .i_b(w_carry_47_13), .i_c(w_carry_47_11), .ow_sum(w_sum_48_15), .ow_carry(w_carry_48_15));
wire w_sum_48_13, w_carry_48_13;
math_adder_full FA_48_13(.i_a(w_carry_47_09), .i_b(w_carry_47_07), .i_c(w_carry_47_05), .ow_sum(w_sum_48_13), .ow_carry(w_carry_48_13));
wire w_sum_48_11, w_carry_48_11;
math_adder_full FA_48_11(.i_a(w_carry_47_03), .i_b(w_sum_48_31), .i_c(w_sum_48_29), .ow_sum(w_sum_48_11), .ow_carry(w_carry_48_11));
wire w_sum_48_09, w_carry_48_09;
math_adder_full FA_48_09(.i_a(w_sum_48_27), .i_b(w_sum_48_25), .i_c(w_sum_48_23), .ow_sum(w_sum_48_09), .ow_carry(w_carry_48_09));
wire w_sum_48_07, w_carry_48_07;
math_adder_full FA_48_07(.i_a(w_sum_48_21), .i_b(w_sum_48_19), .i_c(w_sum_48_17), .ow_sum(w_sum_48_07), .ow_carry(w_carry_48_07));
wire w_sum_48_05, w_carry_48_05;
math_adder_full FA_48_05(.i_a(w_sum_48_15), .i_b(w_sum_48_13), .i_c(w_sum_48_11), .ow_sum(w_sum_48_05), .ow_carry(w_carry_48_05));
wire w_sum_48_03, w_carry_48_03;
math_adder_full FA_48_03(.i_a(w_sum_48_09), .i_b(w_sum_48_07), .i_c(w_sum_48_05), .ow_sum(w_sum_48_03), .ow_carry(w_carry_48_03));
wire w_sum_49_29, w_carry_49_29;
math_adder_full FA_49_29(.i_a(w_pp_18_31), .i_b(w_pp_19_30), .i_c(w_pp_20_29), .ow_sum(w_sum_49_29), .ow_carry(w_carry_49_29));
wire w_sum_49_27, w_carry_49_27;
math_adder_full FA_49_27(.i_a(w_pp_21_28), .i_b(w_pp_22_27), .i_c(w_pp_23_26), .ow_sum(w_sum_49_27), .ow_carry(w_carry_49_27));
wire w_sum_49_25, w_carry_49_25;
math_adder_full FA_49_25(.i_a(w_pp_24_25), .i_b(w_pp_25_24), .i_c(w_pp_26_23), .ow_sum(w_sum_49_25), .ow_carry(w_carry_49_25));
wire w_sum_49_23, w_carry_49_23;
math_adder_full FA_49_23(.i_a(w_pp_27_22), .i_b(w_pp_28_21), .i_c(w_pp_29_20), .ow_sum(w_sum_49_23), .ow_carry(w_carry_49_23));
wire w_sum_49_21, w_carry_49_21;
math_adder_full FA_49_21(.i_a(w_pp_30_19), .i_b(w_pp_31_18), .i_c(w_carry_48_31), .ow_sum(w_sum_49_21), .ow_carry(w_carry_49_21));
wire w_sum_49_19, w_carry_49_19;
math_adder_full FA_49_19(.i_a(w_carry_48_29), .i_b(w_carry_48_27), .i_c(w_carry_48_25), .ow_sum(w_sum_49_19), .ow_carry(w_carry_49_19));
wire w_sum_49_17, w_carry_49_17;
math_adder_full FA_49_17(.i_a(w_carry_48_23), .i_b(w_carry_48_21), .i_c(w_carry_48_19), .ow_sum(w_sum_49_17), .ow_carry(w_carry_49_17));
wire w_sum_49_15, w_carry_49_15;
math_adder_full FA_49_15(.i_a(w_carry_48_17), .i_b(w_carry_48_15), .i_c(w_carry_48_13), .ow_sum(w_sum_49_15), .ow_carry(w_carry_49_15));
wire w_sum_49_13, w_carry_49_13;
math_adder_full FA_49_13(.i_a(w_carry_48_11), .i_b(w_carry_48_09), .i_c(w_carry_48_07), .ow_sum(w_sum_49_13), .ow_carry(w_carry_49_13));
wire w_sum_49_11, w_carry_49_11;
math_adder_full FA_49_11(.i_a(w_carry_48_05), .i_b(w_carry_48_03), .i_c(w_sum_49_29), .ow_sum(w_sum_49_11), .ow_carry(w_carry_49_11));
wire w_sum_49_09, w_carry_49_09;
math_adder_full FA_49_09(.i_a(w_sum_49_27), .i_b(w_sum_49_25), .i_c(w_sum_49_23), .ow_sum(w_sum_49_09), .ow_carry(w_carry_49_09));
wire w_sum_49_07, w_carry_49_07;
math_adder_full FA_49_07(.i_a(w_sum_49_21), .i_b(w_sum_49_19), .i_c(w_sum_49_17), .ow_sum(w_sum_49_07), .ow_carry(w_carry_49_07));
wire w_sum_49_05, w_carry_49_05;
math_adder_full FA_49_05(.i_a(w_sum_49_15), .i_b(w_sum_49_13), .i_c(w_sum_49_11), .ow_sum(w_sum_49_05), .ow_carry(w_carry_49_05));
wire w_sum_49_03, w_carry_49_03;
math_adder_full FA_49_03(.i_a(w_sum_49_09), .i_b(w_sum_49_07), .i_c(w_sum_49_05), .ow_sum(w_sum_49_03), .ow_carry(w_carry_49_03));
wire w_sum_50_27, w_carry_50_27;
math_adder_full FA_50_27(.i_a(w_pp_19_31), .i_b(w_pp_20_30), .i_c(w_pp_21_29), .ow_sum(w_sum_50_27), .ow_carry(w_carry_50_27));
wire w_sum_50_25, w_carry_50_25;
math_adder_full FA_50_25(.i_a(w_pp_22_28), .i_b(w_pp_23_27), .i_c(w_pp_24_26), .ow_sum(w_sum_50_25), .ow_carry(w_carry_50_25));
wire w_sum_50_23, w_carry_50_23;
math_adder_full FA_50_23(.i_a(w_pp_25_25), .i_b(w_pp_26_24), .i_c(w_pp_27_23), .ow_sum(w_sum_50_23), .ow_carry(w_carry_50_23));
wire w_sum_50_21, w_carry_50_21;
math_adder_full FA_50_21(.i_a(w_pp_28_22), .i_b(w_pp_29_21), .i_c(w_pp_30_20), .ow_sum(w_sum_50_21), .ow_carry(w_carry_50_21));
wire w_sum_50_19, w_carry_50_19;
math_adder_full FA_50_19(.i_a(w_pp_31_19), .i_b(w_carry_49_29), .i_c(w_carry_49_27), .ow_sum(w_sum_50_19), .ow_carry(w_carry_50_19));
wire w_sum_50_17, w_carry_50_17;
math_adder_full FA_50_17(.i_a(w_carry_49_25), .i_b(w_carry_49_23), .i_c(w_carry_49_21), .ow_sum(w_sum_50_17), .ow_carry(w_carry_50_17));
wire w_sum_50_15, w_carry_50_15;
math_adder_full FA_50_15(.i_a(w_carry_49_19), .i_b(w_carry_49_17), .i_c(w_carry_49_15), .ow_sum(w_sum_50_15), .ow_carry(w_carry_50_15));
wire w_sum_50_13, w_carry_50_13;
math_adder_full FA_50_13(.i_a(w_carry_49_13), .i_b(w_carry_49_11), .i_c(w_carry_49_09), .ow_sum(w_sum_50_13), .ow_carry(w_carry_50_13));
wire w_sum_50_11, w_carry_50_11;
math_adder_full FA_50_11(.i_a(w_carry_49_07), .i_b(w_carry_49_05), .i_c(w_carry_49_03), .ow_sum(w_sum_50_11), .ow_carry(w_carry_50_11));
wire w_sum_50_09, w_carry_50_09;
math_adder_full FA_50_09(.i_a(w_sum_50_27), .i_b(w_sum_50_25), .i_c(w_sum_50_23), .ow_sum(w_sum_50_09), .ow_carry(w_carry_50_09));
wire w_sum_50_07, w_carry_50_07;
math_adder_full FA_50_07(.i_a(w_sum_50_21), .i_b(w_sum_50_19), .i_c(w_sum_50_17), .ow_sum(w_sum_50_07), .ow_carry(w_carry_50_07));
wire w_sum_50_05, w_carry_50_05;
math_adder_full FA_50_05(.i_a(w_sum_50_15), .i_b(w_sum_50_13), .i_c(w_sum_50_11), .ow_sum(w_sum_50_05), .ow_carry(w_carry_50_05));
wire w_sum_50_03, w_carry_50_03;
math_adder_full FA_50_03(.i_a(w_sum_50_09), .i_b(w_sum_50_07), .i_c(w_sum_50_05), .ow_sum(w_sum_50_03), .ow_carry(w_carry_50_03));
wire w_sum_51_25, w_carry_51_25;
math_adder_full FA_51_25(.i_a(w_pp_20_31), .i_b(w_pp_21_30), .i_c(w_pp_22_29), .ow_sum(w_sum_51_25), .ow_carry(w_carry_51_25));
wire w_sum_51_23, w_carry_51_23;
math_adder_full FA_51_23(.i_a(w_pp_23_28), .i_b(w_pp_24_27), .i_c(w_pp_25_26), .ow_sum(w_sum_51_23), .ow_carry(w_carry_51_23));
wire w_sum_51_21, w_carry_51_21;
math_adder_full FA_51_21(.i_a(w_pp_26_25), .i_b(w_pp_27_24), .i_c(w_pp_28_23), .ow_sum(w_sum_51_21), .ow_carry(w_carry_51_21));
wire w_sum_51_19, w_carry_51_19;
math_adder_full FA_51_19(.i_a(w_pp_29_22), .i_b(w_pp_30_21), .i_c(w_pp_31_20), .ow_sum(w_sum_51_19), .ow_carry(w_carry_51_19));
wire w_sum_51_17, w_carry_51_17;
math_adder_full FA_51_17(.i_a(w_carry_50_27), .i_b(w_carry_50_25), .i_c(w_carry_50_23), .ow_sum(w_sum_51_17), .ow_carry(w_carry_51_17));
wire w_sum_51_15, w_carry_51_15;
math_adder_full FA_51_15(.i_a(w_carry_50_21), .i_b(w_carry_50_19), .i_c(w_carry_50_17), .ow_sum(w_sum_51_15), .ow_carry(w_carry_51_15));
wire w_sum_51_13, w_carry_51_13;
math_adder_full FA_51_13(.i_a(w_carry_50_15), .i_b(w_carry_50_13), .i_c(w_carry_50_11), .ow_sum(w_sum_51_13), .ow_carry(w_carry_51_13));
wire w_sum_51_11, w_carry_51_11;
math_adder_full FA_51_11(.i_a(w_carry_50_09), .i_b(w_carry_50_07), .i_c(w_carry_50_05), .ow_sum(w_sum_51_11), .ow_carry(w_carry_51_11));
wire w_sum_51_09, w_carry_51_09;
math_adder_full FA_51_09(.i_a(w_carry_50_03), .i_b(w_sum_51_25), .i_c(w_sum_51_23), .ow_sum(w_sum_51_09), .ow_carry(w_carry_51_09));
wire w_sum_51_07, w_carry_51_07;
math_adder_full FA_51_07(.i_a(w_sum_51_21), .i_b(w_sum_51_19), .i_c(w_sum_51_17), .ow_sum(w_sum_51_07), .ow_carry(w_carry_51_07));
wire w_sum_51_05, w_carry_51_05;
math_adder_full FA_51_05(.i_a(w_sum_51_15), .i_b(w_sum_51_13), .i_c(w_sum_51_11), .ow_sum(w_sum_51_05), .ow_carry(w_carry_51_05));
wire w_sum_51_03, w_carry_51_03;
math_adder_full FA_51_03(.i_a(w_sum_51_09), .i_b(w_sum_51_07), .i_c(w_sum_51_05), .ow_sum(w_sum_51_03), .ow_carry(w_carry_51_03));
wire w_sum_52_23, w_carry_52_23;
math_adder_full FA_52_23(.i_a(w_pp_21_31), .i_b(w_pp_22_30), .i_c(w_pp_23_29), .ow_sum(w_sum_52_23), .ow_carry(w_carry_52_23));
wire w_sum_52_21, w_carry_52_21;
math_adder_full FA_52_21(.i_a(w_pp_24_28), .i_b(w_pp_25_27), .i_c(w_pp_26_26), .ow_sum(w_sum_52_21), .ow_carry(w_carry_52_21));
wire w_sum_52_19, w_carry_52_19;
math_adder_full FA_52_19(.i_a(w_pp_27_25), .i_b(w_pp_28_24), .i_c(w_pp_29_23), .ow_sum(w_sum_52_19), .ow_carry(w_carry_52_19));
wire w_sum_52_17, w_carry_52_17;
math_adder_full FA_52_17(.i_a(w_pp_30_22), .i_b(w_pp_31_21), .i_c(w_carry_51_25), .ow_sum(w_sum_52_17), .ow_carry(w_carry_52_17));
wire w_sum_52_15, w_carry_52_15;
math_adder_full FA_52_15(.i_a(w_carry_51_23), .i_b(w_carry_51_21), .i_c(w_carry_51_19), .ow_sum(w_sum_52_15), .ow_carry(w_carry_52_15));
wire w_sum_52_13, w_carry_52_13;
math_adder_full FA_52_13(.i_a(w_carry_51_17), .i_b(w_carry_51_15), .i_c(w_carry_51_13), .ow_sum(w_sum_52_13), .ow_carry(w_carry_52_13));
wire w_sum_52_11, w_carry_52_11;
math_adder_full FA_52_11(.i_a(w_carry_51_11), .i_b(w_carry_51_09), .i_c(w_carry_51_07), .ow_sum(w_sum_52_11), .ow_carry(w_carry_52_11));
wire w_sum_52_09, w_carry_52_09;
math_adder_full FA_52_09(.i_a(w_carry_51_05), .i_b(w_carry_51_03), .i_c(w_sum_52_23), .ow_sum(w_sum_52_09), .ow_carry(w_carry_52_09));
wire w_sum_52_07, w_carry_52_07;
math_adder_full FA_52_07(.i_a(w_sum_52_21), .i_b(w_sum_52_19), .i_c(w_sum_52_17), .ow_sum(w_sum_52_07), .ow_carry(w_carry_52_07));
wire w_sum_52_05, w_carry_52_05;
math_adder_full FA_52_05(.i_a(w_sum_52_15), .i_b(w_sum_52_13), .i_c(w_sum_52_11), .ow_sum(w_sum_52_05), .ow_carry(w_carry_52_05));
wire w_sum_52_03, w_carry_52_03;
math_adder_full FA_52_03(.i_a(w_sum_52_09), .i_b(w_sum_52_07), .i_c(w_sum_52_05), .ow_sum(w_sum_52_03), .ow_carry(w_carry_52_03));
wire w_sum_53_21, w_carry_53_21;
math_adder_full FA_53_21(.i_a(w_pp_22_31), .i_b(w_pp_23_30), .i_c(w_pp_24_29), .ow_sum(w_sum_53_21), .ow_carry(w_carry_53_21));
wire w_sum_53_19, w_carry_53_19;
math_adder_full FA_53_19(.i_a(w_pp_25_28), .i_b(w_pp_26_27), .i_c(w_pp_27_26), .ow_sum(w_sum_53_19), .ow_carry(w_carry_53_19));
wire w_sum_53_17, w_carry_53_17;
math_adder_full FA_53_17(.i_a(w_pp_28_25), .i_b(w_pp_29_24), .i_c(w_pp_30_23), .ow_sum(w_sum_53_17), .ow_carry(w_carry_53_17));
wire w_sum_53_15, w_carry_53_15;
math_adder_full FA_53_15(.i_a(w_pp_31_22), .i_b(w_carry_52_23), .i_c(w_carry_52_21), .ow_sum(w_sum_53_15), .ow_carry(w_carry_53_15));
wire w_sum_53_13, w_carry_53_13;
math_adder_full FA_53_13(.i_a(w_carry_52_19), .i_b(w_carry_52_17), .i_c(w_carry_52_15), .ow_sum(w_sum_53_13), .ow_carry(w_carry_53_13));
wire w_sum_53_11, w_carry_53_11;
math_adder_full FA_53_11(.i_a(w_carry_52_13), .i_b(w_carry_52_11), .i_c(w_carry_52_09), .ow_sum(w_sum_53_11), .ow_carry(w_carry_53_11));
wire w_sum_53_09, w_carry_53_09;
math_adder_full FA_53_09(.i_a(w_carry_52_07), .i_b(w_carry_52_05), .i_c(w_carry_52_03), .ow_sum(w_sum_53_09), .ow_carry(w_carry_53_09));
wire w_sum_53_07, w_carry_53_07;
math_adder_full FA_53_07(.i_a(w_sum_53_21), .i_b(w_sum_53_19), .i_c(w_sum_53_17), .ow_sum(w_sum_53_07), .ow_carry(w_carry_53_07));
wire w_sum_53_05, w_carry_53_05;
math_adder_full FA_53_05(.i_a(w_sum_53_15), .i_b(w_sum_53_13), .i_c(w_sum_53_11), .ow_sum(w_sum_53_05), .ow_carry(w_carry_53_05));
wire w_sum_53_03, w_carry_53_03;
math_adder_full FA_53_03(.i_a(w_sum_53_09), .i_b(w_sum_53_07), .i_c(w_sum_53_05), .ow_sum(w_sum_53_03), .ow_carry(w_carry_53_03));
wire w_sum_54_19, w_carry_54_19;
math_adder_full FA_54_19(.i_a(w_pp_23_31), .i_b(w_pp_24_30), .i_c(w_pp_25_29), .ow_sum(w_sum_54_19), .ow_carry(w_carry_54_19));
wire w_sum_54_17, w_carry_54_17;
math_adder_full FA_54_17(.i_a(w_pp_26_28), .i_b(w_pp_27_27), .i_c(w_pp_28_26), .ow_sum(w_sum_54_17), .ow_carry(w_carry_54_17));
wire w_sum_54_15, w_carry_54_15;
math_adder_full FA_54_15(.i_a(w_pp_29_25), .i_b(w_pp_30_24), .i_c(w_pp_31_23), .ow_sum(w_sum_54_15), .ow_carry(w_carry_54_15));
wire w_sum_54_13, w_carry_54_13;
math_adder_full FA_54_13(.i_a(w_carry_53_21), .i_b(w_carry_53_19), .i_c(w_carry_53_17), .ow_sum(w_sum_54_13), .ow_carry(w_carry_54_13));
wire w_sum_54_11, w_carry_54_11;
math_adder_full FA_54_11(.i_a(w_carry_53_15), .i_b(w_carry_53_13), .i_c(w_carry_53_11), .ow_sum(w_sum_54_11), .ow_carry(w_carry_54_11));
wire w_sum_54_09, w_carry_54_09;
math_adder_full FA_54_09(.i_a(w_carry_53_09), .i_b(w_carry_53_07), .i_c(w_carry_53_05), .ow_sum(w_sum_54_09), .ow_carry(w_carry_54_09));
wire w_sum_54_07, w_carry_54_07;
math_adder_full FA_54_07(.i_a(w_carry_53_03), .i_b(w_sum_54_19), .i_c(w_sum_54_17), .ow_sum(w_sum_54_07), .ow_carry(w_carry_54_07));
wire w_sum_54_05, w_carry_54_05;
math_adder_full FA_54_05(.i_a(w_sum_54_15), .i_b(w_sum_54_13), .i_c(w_sum_54_11), .ow_sum(w_sum_54_05), .ow_carry(w_carry_54_05));
wire w_sum_54_03, w_carry_54_03;
math_adder_full FA_54_03(.i_a(w_sum_54_09), .i_b(w_sum_54_07), .i_c(w_sum_54_05), .ow_sum(w_sum_54_03), .ow_carry(w_carry_54_03));
wire w_sum_55_17, w_carry_55_17;
math_adder_full FA_55_17(.i_a(w_pp_24_31), .i_b(w_pp_25_30), .i_c(w_pp_26_29), .ow_sum(w_sum_55_17), .ow_carry(w_carry_55_17));
wire w_sum_55_15, w_carry_55_15;
math_adder_full FA_55_15(.i_a(w_pp_27_28), .i_b(w_pp_28_27), .i_c(w_pp_29_26), .ow_sum(w_sum_55_15), .ow_carry(w_carry_55_15));
wire w_sum_55_13, w_carry_55_13;
math_adder_full FA_55_13(.i_a(w_pp_30_25), .i_b(w_pp_31_24), .i_c(w_carry_54_19), .ow_sum(w_sum_55_13), .ow_carry(w_carry_55_13));
wire w_sum_55_11, w_carry_55_11;
math_adder_full FA_55_11(.i_a(w_carry_54_17), .i_b(w_carry_54_15), .i_c(w_carry_54_13), .ow_sum(w_sum_55_11), .ow_carry(w_carry_55_11));
wire w_sum_55_09, w_carry_55_09;
math_adder_full FA_55_09(.i_a(w_carry_54_11), .i_b(w_carry_54_09), .i_c(w_carry_54_07), .ow_sum(w_sum_55_09), .ow_carry(w_carry_55_09));
wire w_sum_55_07, w_carry_55_07;
math_adder_full FA_55_07(.i_a(w_carry_54_05), .i_b(w_carry_54_03), .i_c(w_sum_55_17), .ow_sum(w_sum_55_07), .ow_carry(w_carry_55_07));
wire w_sum_55_05, w_carry_55_05;
math_adder_full FA_55_05(.i_a(w_sum_55_15), .i_b(w_sum_55_13), .i_c(w_sum_55_11), .ow_sum(w_sum_55_05), .ow_carry(w_carry_55_05));
wire w_sum_55_03, w_carry_55_03;
math_adder_full FA_55_03(.i_a(w_sum_55_09), .i_b(w_sum_55_07), .i_c(w_sum_55_05), .ow_sum(w_sum_55_03), .ow_carry(w_carry_55_03));
wire w_sum_56_15, w_carry_56_15;
math_adder_full FA_56_15(.i_a(w_pp_25_31), .i_b(w_pp_26_30), .i_c(w_pp_27_29), .ow_sum(w_sum_56_15), .ow_carry(w_carry_56_15));
wire w_sum_56_13, w_carry_56_13;
math_adder_full FA_56_13(.i_a(w_pp_28_28), .i_b(w_pp_29_27), .i_c(w_pp_30_26), .ow_sum(w_sum_56_13), .ow_carry(w_carry_56_13));
wire w_sum_56_11, w_carry_56_11;
math_adder_full FA_56_11(.i_a(w_pp_31_25), .i_b(w_carry_55_17), .i_c(w_carry_55_15), .ow_sum(w_sum_56_11), .ow_carry(w_carry_56_11));
wire w_sum_56_09, w_carry_56_09;
math_adder_full FA_56_09(.i_a(w_carry_55_13), .i_b(w_carry_55_11), .i_c(w_carry_55_09), .ow_sum(w_sum_56_09), .ow_carry(w_carry_56_09));
wire w_sum_56_07, w_carry_56_07;
math_adder_full FA_56_07(.i_a(w_carry_55_07), .i_b(w_carry_55_05), .i_c(w_carry_55_03), .ow_sum(w_sum_56_07), .ow_carry(w_carry_56_07));
wire w_sum_56_05, w_carry_56_05;
math_adder_full FA_56_05(.i_a(w_sum_56_15), .i_b(w_sum_56_13), .i_c(w_sum_56_11), .ow_sum(w_sum_56_05), .ow_carry(w_carry_56_05));
wire w_sum_56_03, w_carry_56_03;
math_adder_full FA_56_03(.i_a(w_sum_56_09), .i_b(w_sum_56_07), .i_c(w_sum_56_05), .ow_sum(w_sum_56_03), .ow_carry(w_carry_56_03));
wire w_sum_57_13, w_carry_57_13;
math_adder_full FA_57_13(.i_a(w_pp_26_31), .i_b(w_pp_27_30), .i_c(w_pp_28_29), .ow_sum(w_sum_57_13), .ow_carry(w_carry_57_13));
wire w_sum_57_11, w_carry_57_11;
math_adder_full FA_57_11(.i_a(w_pp_29_28), .i_b(w_pp_30_27), .i_c(w_pp_31_26), .ow_sum(w_sum_57_11), .ow_carry(w_carry_57_11));
wire w_sum_57_09, w_carry_57_09;
math_adder_full FA_57_09(.i_a(w_carry_56_15), .i_b(w_carry_56_13), .i_c(w_carry_56_11), .ow_sum(w_sum_57_09), .ow_carry(w_carry_57_09));
wire w_sum_57_07, w_carry_57_07;
math_adder_full FA_57_07(.i_a(w_carry_56_09), .i_b(w_carry_56_07), .i_c(w_carry_56_05), .ow_sum(w_sum_57_07), .ow_carry(w_carry_57_07));
wire w_sum_57_05, w_carry_57_05;
math_adder_full FA_57_05(.i_a(w_carry_56_03), .i_b(w_sum_57_13), .i_c(w_sum_57_11), .ow_sum(w_sum_57_05), .ow_carry(w_carry_57_05));
wire w_sum_57_03, w_carry_57_03;
math_adder_full FA_57_03(.i_a(w_sum_57_09), .i_b(w_sum_57_07), .i_c(w_sum_57_05), .ow_sum(w_sum_57_03), .ow_carry(w_carry_57_03));
wire w_sum_58_11, w_carry_58_11;
math_adder_full FA_58_11(.i_a(w_pp_27_31), .i_b(w_pp_28_30), .i_c(w_pp_29_29), .ow_sum(w_sum_58_11), .ow_carry(w_carry_58_11));
wire w_sum_58_09, w_carry_58_09;
math_adder_full FA_58_09(.i_a(w_pp_30_28), .i_b(w_pp_31_27), .i_c(w_carry_57_13), .ow_sum(w_sum_58_09), .ow_carry(w_carry_58_09));
wire w_sum_58_07, w_carry_58_07;
math_adder_full FA_58_07(.i_a(w_carry_57_11), .i_b(w_carry_57_09), .i_c(w_carry_57_07), .ow_sum(w_sum_58_07), .ow_carry(w_carry_58_07));
wire w_sum_58_05, w_carry_58_05;
math_adder_full FA_58_05(.i_a(w_carry_57_05), .i_b(w_carry_57_03), .i_c(w_sum_58_11), .ow_sum(w_sum_58_05), .ow_carry(w_carry_58_05));
wire w_sum_58_03, w_carry_58_03;
math_adder_full FA_58_03(.i_a(w_sum_58_09), .i_b(w_sum_58_07), .i_c(w_sum_58_05), .ow_sum(w_sum_58_03), .ow_carry(w_carry_58_03));
wire w_sum_59_09, w_carry_59_09;
math_adder_full FA_59_09(.i_a(w_pp_28_31), .i_b(w_pp_29_30), .i_c(w_pp_30_29), .ow_sum(w_sum_59_09), .ow_carry(w_carry_59_09));
wire w_sum_59_07, w_carry_59_07;
math_adder_full FA_59_07(.i_a(w_pp_31_28), .i_b(w_carry_58_11), .i_c(w_carry_58_09), .ow_sum(w_sum_59_07), .ow_carry(w_carry_59_07));
wire w_sum_59_05, w_carry_59_05;
math_adder_full FA_59_05(.i_a(w_carry_58_07), .i_b(w_carry_58_05), .i_c(w_carry_58_03), .ow_sum(w_sum_59_05), .ow_carry(w_carry_59_05));
wire w_sum_59_03, w_carry_59_03;
math_adder_full FA_59_03(.i_a(w_sum_59_09), .i_b(w_sum_59_07), .i_c(w_sum_59_05), .ow_sum(w_sum_59_03), .ow_carry(w_carry_59_03));
wire w_sum_60_07, w_carry_60_07;
math_adder_full FA_60_07(.i_a(w_pp_29_31), .i_b(w_pp_30_30), .i_c(w_pp_31_29), .ow_sum(w_sum_60_07), .ow_carry(w_carry_60_07));
wire w_sum_60_05, w_carry_60_05;
math_adder_full FA_60_05(.i_a(w_carry_59_09), .i_b(w_carry_59_07), .i_c(w_carry_59_05), .ow_sum(w_sum_60_05), .ow_carry(w_carry_60_05));
wire w_sum_60_03, w_carry_60_03;
math_adder_full FA_60_03(.i_a(w_carry_59_03), .i_b(w_sum_60_07), .i_c(w_sum_60_05), .ow_sum(w_sum_60_03), .ow_carry(w_carry_60_03));
wire w_sum_61_05, w_carry_61_05;
math_adder_full FA_61_05(.i_a(w_pp_30_31), .i_b(w_pp_31_30), .i_c(w_carry_60_07), .ow_sum(w_sum_61_05), .ow_carry(w_carry_61_05));
wire w_sum_61_03, w_carry_61_03;
math_adder_full FA_61_03(.i_a(w_carry_60_05), .i_b(w_carry_60_03), .i_c(w_sum_61_05), .ow_sum(w_sum_61_03), .ow_carry(w_carry_61_03));
wire w_sum_62_03, w_carry_62_03;
math_adder_full FA_62_03(.i_a(w_pp_31_31), .i_b(w_carry_61_05), .i_c(w_carry_61_03), .ow_sum(w_sum_62_03), .ow_carry(w_carry_62_03));

// Final addition stage
wire of_sum_00, of_carry_00;
assign of_sum_00 = w_pp_00_00;
assign of_carry_00 = 1'b0;
wire of_sum_01, of_carry_01;
assign of_sum_01 = w_sum_01_02;
assign of_carry_01 = 1'b0;
wire of_sum_02, of_carry_02;
assign of_sum_02 = w_sum_02_02;
assign of_carry_02 = 1'b0;
wire of_sum_03, of_carry_03;
assign of_sum_03 = w_sum_03_02;
assign of_carry_03 = 1'b0;
wire of_sum_04, of_carry_04;
assign of_sum_04 = w_sum_04_02;
assign of_carry_04 = 1'b0;
wire of_sum_05, of_carry_05;
assign of_sum_05 = w_sum_05_02;
assign of_carry_05 = 1'b0;
wire of_sum_06, of_carry_06;
assign of_sum_06 = w_sum_06_02;
assign of_carry_06 = 1'b0;
wire of_sum_07, of_carry_07;
assign of_sum_07 = w_sum_07_02;
assign of_carry_07 = 1'b0;
wire of_sum_08, of_carry_08;
assign of_sum_08 = w_sum_08_02;
assign of_carry_08 = 1'b0;
wire of_sum_09, of_carry_09;
assign of_sum_09 = w_sum_09_02;
assign of_carry_09 = 1'b0;
wire of_sum_10, of_carry_10;
assign of_sum_10 = w_sum_10_02;
assign of_carry_10 = 1'b0;
wire of_sum_11, of_carry_11;
assign of_sum_11 = w_sum_11_02;
assign of_carry_11 = 1'b0;
wire of_sum_12, of_carry_12;
assign of_sum_12 = w_sum_12_02;
assign of_carry_12 = 1'b0;
wire of_sum_13, of_carry_13;
assign of_sum_13 = w_sum_13_02;
assign of_carry_13 = 1'b0;
wire of_sum_14, of_carry_14;
assign of_sum_14 = w_sum_14_02;
assign of_carry_14 = 1'b0;
wire of_sum_15, of_carry_15;
assign of_sum_15 = w_sum_15_02;
assign of_carry_15 = 1'b0;
wire of_sum_16, of_carry_16;
assign of_sum_16 = w_sum_16_02;
assign of_carry_16 = 1'b0;
wire of_sum_17, of_carry_17;
assign of_sum_17 = w_sum_17_02;
assign of_carry_17 = 1'b0;
wire of_sum_18, of_carry_18;
assign of_sum_18 = w_sum_18_02;
assign of_carry_18 = 1'b0;
wire of_sum_19, of_carry_19;
assign of_sum_19 = w_sum_19_02;
assign of_carry_19 = 1'b0;
wire of_sum_20, of_carry_20;
assign of_sum_20 = w_sum_20_02;
assign of_carry_20 = 1'b0;
wire of_sum_21, of_carry_21;
assign of_sum_21 = w_sum_21_02;
assign of_carry_21 = 1'b0;
wire of_sum_22, of_carry_22;
assign of_sum_22 = w_sum_22_02;
assign of_carry_22 = 1'b0;
wire of_sum_23, of_carry_23;
assign of_sum_23 = w_sum_23_02;
assign of_carry_23 = 1'b0;
wire of_sum_24, of_carry_24;
assign of_sum_24 = w_sum_24_02;
assign of_carry_24 = 1'b0;
wire of_sum_25, of_carry_25;
assign of_sum_25 = w_sum_25_02;
assign of_carry_25 = 1'b0;
wire of_sum_26, of_carry_26;
assign of_sum_26 = w_sum_26_02;
assign of_carry_26 = 1'b0;
wire of_sum_27, of_carry_27;
assign of_sum_27 = w_sum_27_02;
assign of_carry_27 = 1'b0;
wire of_sum_28, of_carry_28;
assign of_sum_28 = w_sum_28_02;
assign of_carry_28 = 1'b0;
wire of_sum_29, of_carry_29;
assign of_sum_29 = w_sum_29_02;
assign of_carry_29 = 1'b0;
wire of_sum_30, of_carry_30;
assign of_sum_30 = w_sum_30_02;
assign of_carry_30 = 1'b0;
wire of_sum_31, of_carry_31;
assign of_sum_31 = w_sum_31_02;
assign of_carry_31 = 1'b0;
wire of_sum_32, of_carry_32;
assign of_sum_32 = w_sum_32_02;
assign of_carry_32 = 1'b0;
wire of_sum_33, of_carry_33;
assign of_sum_33 = w_sum_33_03;
assign of_carry_33 = 1'b0;
wire of_sum_34, of_carry_34;
assign of_sum_34 = w_sum_34_03;
assign of_carry_34 = 1'b0;
wire of_sum_35, of_carry_35;
assign of_sum_35 = w_sum_35_03;
assign of_carry_35 = 1'b0;
wire of_sum_36, of_carry_36;
assign of_sum_36 = w_sum_36_03;
assign of_carry_36 = 1'b0;
wire of_sum_37, of_carry_37;
assign of_sum_37 = w_sum_37_03;
assign of_carry_37 = 1'b0;
wire of_sum_38, of_carry_38;
assign of_sum_38 = w_sum_38_03;
assign of_carry_38 = 1'b0;
wire of_sum_39, of_carry_39;
assign of_sum_39 = w_sum_39_03;
assign of_carry_39 = 1'b0;
wire of_sum_40, of_carry_40;
assign of_sum_40 = w_sum_40_03;
assign of_carry_40 = 1'b0;
wire of_sum_41, of_carry_41;
assign of_sum_41 = w_sum_41_03;
assign of_carry_41 = 1'b0;
wire of_sum_42, of_carry_42;
assign of_sum_42 = w_sum_42_03;
assign of_carry_42 = 1'b0;
wire of_sum_43, of_carry_43;
assign of_sum_43 = w_sum_43_03;
assign of_carry_43 = 1'b0;
wire of_sum_44, of_carry_44;
assign of_sum_44 = w_sum_44_03;
assign of_carry_44 = 1'b0;
wire of_sum_45, of_carry_45;
assign of_sum_45 = w_sum_45_03;
assign of_carry_45 = 1'b0;
wire of_sum_46, of_carry_46;
assign of_sum_46 = w_sum_46_03;
assign of_carry_46 = 1'b0;
wire of_sum_47, of_carry_47;
assign of_sum_47 = w_sum_47_03;
assign of_carry_47 = 1'b0;
wire of_sum_48, of_carry_48;
assign of_sum_48 = w_sum_48_03;
assign of_carry_48 = 1'b0;
wire of_sum_49, of_carry_49;
assign of_sum_49 = w_sum_49_03;
assign of_carry_49 = 1'b0;
wire of_sum_50, of_carry_50;
assign of_sum_50 = w_sum_50_03;
assign of_carry_50 = 1'b0;
wire of_sum_51, of_carry_51;
assign of_sum_51 = w_sum_51_03;
assign of_carry_51 = 1'b0;
wire of_sum_52, of_carry_52;
assign of_sum_52 = w_sum_52_03;
assign of_carry_52 = 1'b0;
wire of_sum_53, of_carry_53;
assign of_sum_53 = w_sum_53_03;
assign of_carry_53 = 1'b0;
wire of_sum_54, of_carry_54;
assign of_sum_54 = w_sum_54_03;
assign of_carry_54 = 1'b0;
wire of_sum_55, of_carry_55;
assign of_sum_55 = w_sum_55_03;
assign of_carry_55 = 1'b0;
wire of_sum_56, of_carry_56;
assign of_sum_56 = w_sum_56_03;
assign of_carry_56 = 1'b0;
wire of_sum_57, of_carry_57;
assign of_sum_57 = w_sum_57_03;
assign of_carry_57 = 1'b0;
wire of_sum_58, of_carry_58;
assign of_sum_58 = w_sum_58_03;
assign of_carry_58 = 1'b0;
wire of_sum_59, of_carry_59;
assign of_sum_59 = w_sum_59_03;
assign of_carry_59 = 1'b0;
wire of_sum_60, of_carry_60;
assign of_sum_60 = w_sum_60_03;
assign of_carry_60 = 1'b0;
wire of_sum_61, of_carry_61;
assign of_sum_61 = w_sum_61_03;
assign of_carry_61 = 1'b0;
wire of_sum_62, of_carry_62;
assign of_sum_62 = w_sum_62_03;
assign of_carry_62 = 1'b0;
wire of_sum_63, of_carry_63;
assign of_sum_63 = w_carry_62_03;
assign of_carry_63 = 1'b0;

// Final product assignment
assign ow_product[ 0] = of_sum_00;
assign ow_product[ 1] = of_sum_01;
assign ow_product[ 2] = of_sum_02;
assign ow_product[ 3] = of_sum_03;
assign ow_product[ 4] = of_sum_04;
assign ow_product[ 5] = of_sum_05;
assign ow_product[ 6] = of_sum_06;
assign ow_product[ 7] = of_sum_07;
assign ow_product[ 8] = of_sum_08;
assign ow_product[ 9] = of_sum_09;
assign ow_product[10] = of_sum_10;
assign ow_product[11] = of_sum_11;
assign ow_product[12] = of_sum_12;
assign ow_product[13] = of_sum_13;
assign ow_product[14] = of_sum_14;
assign ow_product[15] = of_sum_15;
assign ow_product[16] = of_sum_16;
assign ow_product[17] = of_sum_17;
assign ow_product[18] = of_sum_18;
assign ow_product[19] = of_sum_19;
assign ow_product[20] = of_sum_20;
assign ow_product[21] = of_sum_21;
assign ow_product[22] = of_sum_22;
assign ow_product[23] = of_sum_23;
assign ow_product[24] = of_sum_24;
assign ow_product[25] = of_sum_25;
assign ow_product[26] = of_sum_26;
assign ow_product[27] = of_sum_27;
assign ow_product[28] = of_sum_28;
assign ow_product[29] = of_sum_29;
assign ow_product[30] = of_sum_30;
assign ow_product[31] = of_sum_31;
assign ow_product[32] = of_sum_32;
assign ow_product[33] = of_sum_33;
assign ow_product[34] = of_sum_34;
assign ow_product[35] = of_sum_35;
assign ow_product[36] = of_sum_36;
assign ow_product[37] = of_sum_37;
assign ow_product[38] = of_sum_38;
assign ow_product[39] = of_sum_39;
assign ow_product[40] = of_sum_40;
assign ow_product[41] = of_sum_41;
assign ow_product[42] = of_sum_42;
assign ow_product[43] = of_sum_43;
assign ow_product[44] = of_sum_44;
assign ow_product[45] = of_sum_45;
assign ow_product[46] = of_sum_46;
assign ow_product[47] = of_sum_47;
assign ow_product[48] = of_sum_48;
assign ow_product[49] = of_sum_49;
assign ow_product[50] = of_sum_50;
assign ow_product[51] = of_sum_51;
assign ow_product[52] = of_sum_52;
assign ow_product[53] = of_sum_53;
assign ow_product[54] = of_sum_54;
assign ow_product[55] = of_sum_55;
assign ow_product[56] = of_sum_56;
assign ow_product[57] = of_sum_57;
assign ow_product[58] = of_sum_58;
assign ow_product[59] = of_sum_59;
assign ow_product[60] = of_sum_60;
assign ow_product[61] = of_sum_61;
assign ow_product[62] = of_sum_62;
assign ow_product[63] = of_sum_63;


    // Debug purposes
    // synopsys translate_off
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_wallace_tree_032);
    end
    // synopsys translate_on
        
endmodule : math_multiplier_wallace_tree_032
