`timescale 1ns / 1ps

module math_multiplier_wallace_tree_csa_32 (
    input  [31:0] i_multiplier,
    input  [31:0] i_multiplicand,
    output [63:0] ow_product
);

// Partial products generation
wire w_pp_0_0 = i_multiplier[0] & i_multiplicand[0];
wire w_pp_0_1 = i_multiplier[0] & i_multiplicand[1];
wire w_pp_0_2 = i_multiplier[0] & i_multiplicand[2];
wire w_pp_0_3 = i_multiplier[0] & i_multiplicand[3];
wire w_pp_0_4 = i_multiplier[0] & i_multiplicand[4];
wire w_pp_0_5 = i_multiplier[0] & i_multiplicand[5];
wire w_pp_0_6 = i_multiplier[0] & i_multiplicand[6];
wire w_pp_0_7 = i_multiplier[0] & i_multiplicand[7];
wire w_pp_0_8 = i_multiplier[0] & i_multiplicand[8];
wire w_pp_0_9 = i_multiplier[0] & i_multiplicand[9];
wire w_pp_0_10 = i_multiplier[0] & i_multiplicand[10];
wire w_pp_0_11 = i_multiplier[0] & i_multiplicand[11];
wire w_pp_0_12 = i_multiplier[0] & i_multiplicand[12];
wire w_pp_0_13 = i_multiplier[0] & i_multiplicand[13];
wire w_pp_0_14 = i_multiplier[0] & i_multiplicand[14];
wire w_pp_0_15 = i_multiplier[0] & i_multiplicand[15];
wire w_pp_0_16 = i_multiplier[0] & i_multiplicand[16];
wire w_pp_0_17 = i_multiplier[0] & i_multiplicand[17];
wire w_pp_0_18 = i_multiplier[0] & i_multiplicand[18];
wire w_pp_0_19 = i_multiplier[0] & i_multiplicand[19];
wire w_pp_0_20 = i_multiplier[0] & i_multiplicand[20];
wire w_pp_0_21 = i_multiplier[0] & i_multiplicand[21];
wire w_pp_0_22 = i_multiplier[0] & i_multiplicand[22];
wire w_pp_0_23 = i_multiplier[0] & i_multiplicand[23];
wire w_pp_0_24 = i_multiplier[0] & i_multiplicand[24];
wire w_pp_0_25 = i_multiplier[0] & i_multiplicand[25];
wire w_pp_0_26 = i_multiplier[0] & i_multiplicand[26];
wire w_pp_0_27 = i_multiplier[0] & i_multiplicand[27];
wire w_pp_0_28 = i_multiplier[0] & i_multiplicand[28];
wire w_pp_0_29 = i_multiplier[0] & i_multiplicand[29];
wire w_pp_0_30 = i_multiplier[0] & i_multiplicand[30];
wire w_pp_0_31 = i_multiplier[0] & i_multiplicand[31];
wire w_pp_1_0 = i_multiplier[1] & i_multiplicand[0];
wire w_pp_1_1 = i_multiplier[1] & i_multiplicand[1];
wire w_pp_1_2 = i_multiplier[1] & i_multiplicand[2];
wire w_pp_1_3 = i_multiplier[1] & i_multiplicand[3];
wire w_pp_1_4 = i_multiplier[1] & i_multiplicand[4];
wire w_pp_1_5 = i_multiplier[1] & i_multiplicand[5];
wire w_pp_1_6 = i_multiplier[1] & i_multiplicand[6];
wire w_pp_1_7 = i_multiplier[1] & i_multiplicand[7];
wire w_pp_1_8 = i_multiplier[1] & i_multiplicand[8];
wire w_pp_1_9 = i_multiplier[1] & i_multiplicand[9];
wire w_pp_1_10 = i_multiplier[1] & i_multiplicand[10];
wire w_pp_1_11 = i_multiplier[1] & i_multiplicand[11];
wire w_pp_1_12 = i_multiplier[1] & i_multiplicand[12];
wire w_pp_1_13 = i_multiplier[1] & i_multiplicand[13];
wire w_pp_1_14 = i_multiplier[1] & i_multiplicand[14];
wire w_pp_1_15 = i_multiplier[1] & i_multiplicand[15];
wire w_pp_1_16 = i_multiplier[1] & i_multiplicand[16];
wire w_pp_1_17 = i_multiplier[1] & i_multiplicand[17];
wire w_pp_1_18 = i_multiplier[1] & i_multiplicand[18];
wire w_pp_1_19 = i_multiplier[1] & i_multiplicand[19];
wire w_pp_1_20 = i_multiplier[1] & i_multiplicand[20];
wire w_pp_1_21 = i_multiplier[1] & i_multiplicand[21];
wire w_pp_1_22 = i_multiplier[1] & i_multiplicand[22];
wire w_pp_1_23 = i_multiplier[1] & i_multiplicand[23];
wire w_pp_1_24 = i_multiplier[1] & i_multiplicand[24];
wire w_pp_1_25 = i_multiplier[1] & i_multiplicand[25];
wire w_pp_1_26 = i_multiplier[1] & i_multiplicand[26];
wire w_pp_1_27 = i_multiplier[1] & i_multiplicand[27];
wire w_pp_1_28 = i_multiplier[1] & i_multiplicand[28];
wire w_pp_1_29 = i_multiplier[1] & i_multiplicand[29];
wire w_pp_1_30 = i_multiplier[1] & i_multiplicand[30];
wire w_pp_1_31 = i_multiplier[1] & i_multiplicand[31];
wire w_pp_2_0 = i_multiplier[2] & i_multiplicand[0];
wire w_pp_2_1 = i_multiplier[2] & i_multiplicand[1];
wire w_pp_2_2 = i_multiplier[2] & i_multiplicand[2];
wire w_pp_2_3 = i_multiplier[2] & i_multiplicand[3];
wire w_pp_2_4 = i_multiplier[2] & i_multiplicand[4];
wire w_pp_2_5 = i_multiplier[2] & i_multiplicand[5];
wire w_pp_2_6 = i_multiplier[2] & i_multiplicand[6];
wire w_pp_2_7 = i_multiplier[2] & i_multiplicand[7];
wire w_pp_2_8 = i_multiplier[2] & i_multiplicand[8];
wire w_pp_2_9 = i_multiplier[2] & i_multiplicand[9];
wire w_pp_2_10 = i_multiplier[2] & i_multiplicand[10];
wire w_pp_2_11 = i_multiplier[2] & i_multiplicand[11];
wire w_pp_2_12 = i_multiplier[2] & i_multiplicand[12];
wire w_pp_2_13 = i_multiplier[2] & i_multiplicand[13];
wire w_pp_2_14 = i_multiplier[2] & i_multiplicand[14];
wire w_pp_2_15 = i_multiplier[2] & i_multiplicand[15];
wire w_pp_2_16 = i_multiplier[2] & i_multiplicand[16];
wire w_pp_2_17 = i_multiplier[2] & i_multiplicand[17];
wire w_pp_2_18 = i_multiplier[2] & i_multiplicand[18];
wire w_pp_2_19 = i_multiplier[2] & i_multiplicand[19];
wire w_pp_2_20 = i_multiplier[2] & i_multiplicand[20];
wire w_pp_2_21 = i_multiplier[2] & i_multiplicand[21];
wire w_pp_2_22 = i_multiplier[2] & i_multiplicand[22];
wire w_pp_2_23 = i_multiplier[2] & i_multiplicand[23];
wire w_pp_2_24 = i_multiplier[2] & i_multiplicand[24];
wire w_pp_2_25 = i_multiplier[2] & i_multiplicand[25];
wire w_pp_2_26 = i_multiplier[2] & i_multiplicand[26];
wire w_pp_2_27 = i_multiplier[2] & i_multiplicand[27];
wire w_pp_2_28 = i_multiplier[2] & i_multiplicand[28];
wire w_pp_2_29 = i_multiplier[2] & i_multiplicand[29];
wire w_pp_2_30 = i_multiplier[2] & i_multiplicand[30];
wire w_pp_2_31 = i_multiplier[2] & i_multiplicand[31];
wire w_pp_3_0 = i_multiplier[3] & i_multiplicand[0];
wire w_pp_3_1 = i_multiplier[3] & i_multiplicand[1];
wire w_pp_3_2 = i_multiplier[3] & i_multiplicand[2];
wire w_pp_3_3 = i_multiplier[3] & i_multiplicand[3];
wire w_pp_3_4 = i_multiplier[3] & i_multiplicand[4];
wire w_pp_3_5 = i_multiplier[3] & i_multiplicand[5];
wire w_pp_3_6 = i_multiplier[3] & i_multiplicand[6];
wire w_pp_3_7 = i_multiplier[3] & i_multiplicand[7];
wire w_pp_3_8 = i_multiplier[3] & i_multiplicand[8];
wire w_pp_3_9 = i_multiplier[3] & i_multiplicand[9];
wire w_pp_3_10 = i_multiplier[3] & i_multiplicand[10];
wire w_pp_3_11 = i_multiplier[3] & i_multiplicand[11];
wire w_pp_3_12 = i_multiplier[3] & i_multiplicand[12];
wire w_pp_3_13 = i_multiplier[3] & i_multiplicand[13];
wire w_pp_3_14 = i_multiplier[3] & i_multiplicand[14];
wire w_pp_3_15 = i_multiplier[3] & i_multiplicand[15];
wire w_pp_3_16 = i_multiplier[3] & i_multiplicand[16];
wire w_pp_3_17 = i_multiplier[3] & i_multiplicand[17];
wire w_pp_3_18 = i_multiplier[3] & i_multiplicand[18];
wire w_pp_3_19 = i_multiplier[3] & i_multiplicand[19];
wire w_pp_3_20 = i_multiplier[3] & i_multiplicand[20];
wire w_pp_3_21 = i_multiplier[3] & i_multiplicand[21];
wire w_pp_3_22 = i_multiplier[3] & i_multiplicand[22];
wire w_pp_3_23 = i_multiplier[3] & i_multiplicand[23];
wire w_pp_3_24 = i_multiplier[3] & i_multiplicand[24];
wire w_pp_3_25 = i_multiplier[3] & i_multiplicand[25];
wire w_pp_3_26 = i_multiplier[3] & i_multiplicand[26];
wire w_pp_3_27 = i_multiplier[3] & i_multiplicand[27];
wire w_pp_3_28 = i_multiplier[3] & i_multiplicand[28];
wire w_pp_3_29 = i_multiplier[3] & i_multiplicand[29];
wire w_pp_3_30 = i_multiplier[3] & i_multiplicand[30];
wire w_pp_3_31 = i_multiplier[3] & i_multiplicand[31];
wire w_pp_4_0 = i_multiplier[4] & i_multiplicand[0];
wire w_pp_4_1 = i_multiplier[4] & i_multiplicand[1];
wire w_pp_4_2 = i_multiplier[4] & i_multiplicand[2];
wire w_pp_4_3 = i_multiplier[4] & i_multiplicand[3];
wire w_pp_4_4 = i_multiplier[4] & i_multiplicand[4];
wire w_pp_4_5 = i_multiplier[4] & i_multiplicand[5];
wire w_pp_4_6 = i_multiplier[4] & i_multiplicand[6];
wire w_pp_4_7 = i_multiplier[4] & i_multiplicand[7];
wire w_pp_4_8 = i_multiplier[4] & i_multiplicand[8];
wire w_pp_4_9 = i_multiplier[4] & i_multiplicand[9];
wire w_pp_4_10 = i_multiplier[4] & i_multiplicand[10];
wire w_pp_4_11 = i_multiplier[4] & i_multiplicand[11];
wire w_pp_4_12 = i_multiplier[4] & i_multiplicand[12];
wire w_pp_4_13 = i_multiplier[4] & i_multiplicand[13];
wire w_pp_4_14 = i_multiplier[4] & i_multiplicand[14];
wire w_pp_4_15 = i_multiplier[4] & i_multiplicand[15];
wire w_pp_4_16 = i_multiplier[4] & i_multiplicand[16];
wire w_pp_4_17 = i_multiplier[4] & i_multiplicand[17];
wire w_pp_4_18 = i_multiplier[4] & i_multiplicand[18];
wire w_pp_4_19 = i_multiplier[4] & i_multiplicand[19];
wire w_pp_4_20 = i_multiplier[4] & i_multiplicand[20];
wire w_pp_4_21 = i_multiplier[4] & i_multiplicand[21];
wire w_pp_4_22 = i_multiplier[4] & i_multiplicand[22];
wire w_pp_4_23 = i_multiplier[4] & i_multiplicand[23];
wire w_pp_4_24 = i_multiplier[4] & i_multiplicand[24];
wire w_pp_4_25 = i_multiplier[4] & i_multiplicand[25];
wire w_pp_4_26 = i_multiplier[4] & i_multiplicand[26];
wire w_pp_4_27 = i_multiplier[4] & i_multiplicand[27];
wire w_pp_4_28 = i_multiplier[4] & i_multiplicand[28];
wire w_pp_4_29 = i_multiplier[4] & i_multiplicand[29];
wire w_pp_4_30 = i_multiplier[4] & i_multiplicand[30];
wire w_pp_4_31 = i_multiplier[4] & i_multiplicand[31];
wire w_pp_5_0 = i_multiplier[5] & i_multiplicand[0];
wire w_pp_5_1 = i_multiplier[5] & i_multiplicand[1];
wire w_pp_5_2 = i_multiplier[5] & i_multiplicand[2];
wire w_pp_5_3 = i_multiplier[5] & i_multiplicand[3];
wire w_pp_5_4 = i_multiplier[5] & i_multiplicand[4];
wire w_pp_5_5 = i_multiplier[5] & i_multiplicand[5];
wire w_pp_5_6 = i_multiplier[5] & i_multiplicand[6];
wire w_pp_5_7 = i_multiplier[5] & i_multiplicand[7];
wire w_pp_5_8 = i_multiplier[5] & i_multiplicand[8];
wire w_pp_5_9 = i_multiplier[5] & i_multiplicand[9];
wire w_pp_5_10 = i_multiplier[5] & i_multiplicand[10];
wire w_pp_5_11 = i_multiplier[5] & i_multiplicand[11];
wire w_pp_5_12 = i_multiplier[5] & i_multiplicand[12];
wire w_pp_5_13 = i_multiplier[5] & i_multiplicand[13];
wire w_pp_5_14 = i_multiplier[5] & i_multiplicand[14];
wire w_pp_5_15 = i_multiplier[5] & i_multiplicand[15];
wire w_pp_5_16 = i_multiplier[5] & i_multiplicand[16];
wire w_pp_5_17 = i_multiplier[5] & i_multiplicand[17];
wire w_pp_5_18 = i_multiplier[5] & i_multiplicand[18];
wire w_pp_5_19 = i_multiplier[5] & i_multiplicand[19];
wire w_pp_5_20 = i_multiplier[5] & i_multiplicand[20];
wire w_pp_5_21 = i_multiplier[5] & i_multiplicand[21];
wire w_pp_5_22 = i_multiplier[5] & i_multiplicand[22];
wire w_pp_5_23 = i_multiplier[5] & i_multiplicand[23];
wire w_pp_5_24 = i_multiplier[5] & i_multiplicand[24];
wire w_pp_5_25 = i_multiplier[5] & i_multiplicand[25];
wire w_pp_5_26 = i_multiplier[5] & i_multiplicand[26];
wire w_pp_5_27 = i_multiplier[5] & i_multiplicand[27];
wire w_pp_5_28 = i_multiplier[5] & i_multiplicand[28];
wire w_pp_5_29 = i_multiplier[5] & i_multiplicand[29];
wire w_pp_5_30 = i_multiplier[5] & i_multiplicand[30];
wire w_pp_5_31 = i_multiplier[5] & i_multiplicand[31];
wire w_pp_6_0 = i_multiplier[6] & i_multiplicand[0];
wire w_pp_6_1 = i_multiplier[6] & i_multiplicand[1];
wire w_pp_6_2 = i_multiplier[6] & i_multiplicand[2];
wire w_pp_6_3 = i_multiplier[6] & i_multiplicand[3];
wire w_pp_6_4 = i_multiplier[6] & i_multiplicand[4];
wire w_pp_6_5 = i_multiplier[6] & i_multiplicand[5];
wire w_pp_6_6 = i_multiplier[6] & i_multiplicand[6];
wire w_pp_6_7 = i_multiplier[6] & i_multiplicand[7];
wire w_pp_6_8 = i_multiplier[6] & i_multiplicand[8];
wire w_pp_6_9 = i_multiplier[6] & i_multiplicand[9];
wire w_pp_6_10 = i_multiplier[6] & i_multiplicand[10];
wire w_pp_6_11 = i_multiplier[6] & i_multiplicand[11];
wire w_pp_6_12 = i_multiplier[6] & i_multiplicand[12];
wire w_pp_6_13 = i_multiplier[6] & i_multiplicand[13];
wire w_pp_6_14 = i_multiplier[6] & i_multiplicand[14];
wire w_pp_6_15 = i_multiplier[6] & i_multiplicand[15];
wire w_pp_6_16 = i_multiplier[6] & i_multiplicand[16];
wire w_pp_6_17 = i_multiplier[6] & i_multiplicand[17];
wire w_pp_6_18 = i_multiplier[6] & i_multiplicand[18];
wire w_pp_6_19 = i_multiplier[6] & i_multiplicand[19];
wire w_pp_6_20 = i_multiplier[6] & i_multiplicand[20];
wire w_pp_6_21 = i_multiplier[6] & i_multiplicand[21];
wire w_pp_6_22 = i_multiplier[6] & i_multiplicand[22];
wire w_pp_6_23 = i_multiplier[6] & i_multiplicand[23];
wire w_pp_6_24 = i_multiplier[6] & i_multiplicand[24];
wire w_pp_6_25 = i_multiplier[6] & i_multiplicand[25];
wire w_pp_6_26 = i_multiplier[6] & i_multiplicand[26];
wire w_pp_6_27 = i_multiplier[6] & i_multiplicand[27];
wire w_pp_6_28 = i_multiplier[6] & i_multiplicand[28];
wire w_pp_6_29 = i_multiplier[6] & i_multiplicand[29];
wire w_pp_6_30 = i_multiplier[6] & i_multiplicand[30];
wire w_pp_6_31 = i_multiplier[6] & i_multiplicand[31];
wire w_pp_7_0 = i_multiplier[7] & i_multiplicand[0];
wire w_pp_7_1 = i_multiplier[7] & i_multiplicand[1];
wire w_pp_7_2 = i_multiplier[7] & i_multiplicand[2];
wire w_pp_7_3 = i_multiplier[7] & i_multiplicand[3];
wire w_pp_7_4 = i_multiplier[7] & i_multiplicand[4];
wire w_pp_7_5 = i_multiplier[7] & i_multiplicand[5];
wire w_pp_7_6 = i_multiplier[7] & i_multiplicand[6];
wire w_pp_7_7 = i_multiplier[7] & i_multiplicand[7];
wire w_pp_7_8 = i_multiplier[7] & i_multiplicand[8];
wire w_pp_7_9 = i_multiplier[7] & i_multiplicand[9];
wire w_pp_7_10 = i_multiplier[7] & i_multiplicand[10];
wire w_pp_7_11 = i_multiplier[7] & i_multiplicand[11];
wire w_pp_7_12 = i_multiplier[7] & i_multiplicand[12];
wire w_pp_7_13 = i_multiplier[7] & i_multiplicand[13];
wire w_pp_7_14 = i_multiplier[7] & i_multiplicand[14];
wire w_pp_7_15 = i_multiplier[7] & i_multiplicand[15];
wire w_pp_7_16 = i_multiplier[7] & i_multiplicand[16];
wire w_pp_7_17 = i_multiplier[7] & i_multiplicand[17];
wire w_pp_7_18 = i_multiplier[7] & i_multiplicand[18];
wire w_pp_7_19 = i_multiplier[7] & i_multiplicand[19];
wire w_pp_7_20 = i_multiplier[7] & i_multiplicand[20];
wire w_pp_7_21 = i_multiplier[7] & i_multiplicand[21];
wire w_pp_7_22 = i_multiplier[7] & i_multiplicand[22];
wire w_pp_7_23 = i_multiplier[7] & i_multiplicand[23];
wire w_pp_7_24 = i_multiplier[7] & i_multiplicand[24];
wire w_pp_7_25 = i_multiplier[7] & i_multiplicand[25];
wire w_pp_7_26 = i_multiplier[7] & i_multiplicand[26];
wire w_pp_7_27 = i_multiplier[7] & i_multiplicand[27];
wire w_pp_7_28 = i_multiplier[7] & i_multiplicand[28];
wire w_pp_7_29 = i_multiplier[7] & i_multiplicand[29];
wire w_pp_7_30 = i_multiplier[7] & i_multiplicand[30];
wire w_pp_7_31 = i_multiplier[7] & i_multiplicand[31];
wire w_pp_8_0 = i_multiplier[8] & i_multiplicand[0];
wire w_pp_8_1 = i_multiplier[8] & i_multiplicand[1];
wire w_pp_8_2 = i_multiplier[8] & i_multiplicand[2];
wire w_pp_8_3 = i_multiplier[8] & i_multiplicand[3];
wire w_pp_8_4 = i_multiplier[8] & i_multiplicand[4];
wire w_pp_8_5 = i_multiplier[8] & i_multiplicand[5];
wire w_pp_8_6 = i_multiplier[8] & i_multiplicand[6];
wire w_pp_8_7 = i_multiplier[8] & i_multiplicand[7];
wire w_pp_8_8 = i_multiplier[8] & i_multiplicand[8];
wire w_pp_8_9 = i_multiplier[8] & i_multiplicand[9];
wire w_pp_8_10 = i_multiplier[8] & i_multiplicand[10];
wire w_pp_8_11 = i_multiplier[8] & i_multiplicand[11];
wire w_pp_8_12 = i_multiplier[8] & i_multiplicand[12];
wire w_pp_8_13 = i_multiplier[8] & i_multiplicand[13];
wire w_pp_8_14 = i_multiplier[8] & i_multiplicand[14];
wire w_pp_8_15 = i_multiplier[8] & i_multiplicand[15];
wire w_pp_8_16 = i_multiplier[8] & i_multiplicand[16];
wire w_pp_8_17 = i_multiplier[8] & i_multiplicand[17];
wire w_pp_8_18 = i_multiplier[8] & i_multiplicand[18];
wire w_pp_8_19 = i_multiplier[8] & i_multiplicand[19];
wire w_pp_8_20 = i_multiplier[8] & i_multiplicand[20];
wire w_pp_8_21 = i_multiplier[8] & i_multiplicand[21];
wire w_pp_8_22 = i_multiplier[8] & i_multiplicand[22];
wire w_pp_8_23 = i_multiplier[8] & i_multiplicand[23];
wire w_pp_8_24 = i_multiplier[8] & i_multiplicand[24];
wire w_pp_8_25 = i_multiplier[8] & i_multiplicand[25];
wire w_pp_8_26 = i_multiplier[8] & i_multiplicand[26];
wire w_pp_8_27 = i_multiplier[8] & i_multiplicand[27];
wire w_pp_8_28 = i_multiplier[8] & i_multiplicand[28];
wire w_pp_8_29 = i_multiplier[8] & i_multiplicand[29];
wire w_pp_8_30 = i_multiplier[8] & i_multiplicand[30];
wire w_pp_8_31 = i_multiplier[8] & i_multiplicand[31];
wire w_pp_9_0 = i_multiplier[9] & i_multiplicand[0];
wire w_pp_9_1 = i_multiplier[9] & i_multiplicand[1];
wire w_pp_9_2 = i_multiplier[9] & i_multiplicand[2];
wire w_pp_9_3 = i_multiplier[9] & i_multiplicand[3];
wire w_pp_9_4 = i_multiplier[9] & i_multiplicand[4];
wire w_pp_9_5 = i_multiplier[9] & i_multiplicand[5];
wire w_pp_9_6 = i_multiplier[9] & i_multiplicand[6];
wire w_pp_9_7 = i_multiplier[9] & i_multiplicand[7];
wire w_pp_9_8 = i_multiplier[9] & i_multiplicand[8];
wire w_pp_9_9 = i_multiplier[9] & i_multiplicand[9];
wire w_pp_9_10 = i_multiplier[9] & i_multiplicand[10];
wire w_pp_9_11 = i_multiplier[9] & i_multiplicand[11];
wire w_pp_9_12 = i_multiplier[9] & i_multiplicand[12];
wire w_pp_9_13 = i_multiplier[9] & i_multiplicand[13];
wire w_pp_9_14 = i_multiplier[9] & i_multiplicand[14];
wire w_pp_9_15 = i_multiplier[9] & i_multiplicand[15];
wire w_pp_9_16 = i_multiplier[9] & i_multiplicand[16];
wire w_pp_9_17 = i_multiplier[9] & i_multiplicand[17];
wire w_pp_9_18 = i_multiplier[9] & i_multiplicand[18];
wire w_pp_9_19 = i_multiplier[9] & i_multiplicand[19];
wire w_pp_9_20 = i_multiplier[9] & i_multiplicand[20];
wire w_pp_9_21 = i_multiplier[9] & i_multiplicand[21];
wire w_pp_9_22 = i_multiplier[9] & i_multiplicand[22];
wire w_pp_9_23 = i_multiplier[9] & i_multiplicand[23];
wire w_pp_9_24 = i_multiplier[9] & i_multiplicand[24];
wire w_pp_9_25 = i_multiplier[9] & i_multiplicand[25];
wire w_pp_9_26 = i_multiplier[9] & i_multiplicand[26];
wire w_pp_9_27 = i_multiplier[9] & i_multiplicand[27];
wire w_pp_9_28 = i_multiplier[9] & i_multiplicand[28];
wire w_pp_9_29 = i_multiplier[9] & i_multiplicand[29];
wire w_pp_9_30 = i_multiplier[9] & i_multiplicand[30];
wire w_pp_9_31 = i_multiplier[9] & i_multiplicand[31];
wire w_pp_10_0 = i_multiplier[10] & i_multiplicand[0];
wire w_pp_10_1 = i_multiplier[10] & i_multiplicand[1];
wire w_pp_10_2 = i_multiplier[10] & i_multiplicand[2];
wire w_pp_10_3 = i_multiplier[10] & i_multiplicand[3];
wire w_pp_10_4 = i_multiplier[10] & i_multiplicand[4];
wire w_pp_10_5 = i_multiplier[10] & i_multiplicand[5];
wire w_pp_10_6 = i_multiplier[10] & i_multiplicand[6];
wire w_pp_10_7 = i_multiplier[10] & i_multiplicand[7];
wire w_pp_10_8 = i_multiplier[10] & i_multiplicand[8];
wire w_pp_10_9 = i_multiplier[10] & i_multiplicand[9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_10_16 = i_multiplier[10] & i_multiplicand[16];
wire w_pp_10_17 = i_multiplier[10] & i_multiplicand[17];
wire w_pp_10_18 = i_multiplier[10] & i_multiplicand[18];
wire w_pp_10_19 = i_multiplier[10] & i_multiplicand[19];
wire w_pp_10_20 = i_multiplier[10] & i_multiplicand[20];
wire w_pp_10_21 = i_multiplier[10] & i_multiplicand[21];
wire w_pp_10_22 = i_multiplier[10] & i_multiplicand[22];
wire w_pp_10_23 = i_multiplier[10] & i_multiplicand[23];
wire w_pp_10_24 = i_multiplier[10] & i_multiplicand[24];
wire w_pp_10_25 = i_multiplier[10] & i_multiplicand[25];
wire w_pp_10_26 = i_multiplier[10] & i_multiplicand[26];
wire w_pp_10_27 = i_multiplier[10] & i_multiplicand[27];
wire w_pp_10_28 = i_multiplier[10] & i_multiplicand[28];
wire w_pp_10_29 = i_multiplier[10] & i_multiplicand[29];
wire w_pp_10_30 = i_multiplier[10] & i_multiplicand[30];
wire w_pp_10_31 = i_multiplier[10] & i_multiplicand[31];
wire w_pp_11_0 = i_multiplier[11] & i_multiplicand[0];
wire w_pp_11_1 = i_multiplier[11] & i_multiplicand[1];
wire w_pp_11_2 = i_multiplier[11] & i_multiplicand[2];
wire w_pp_11_3 = i_multiplier[11] & i_multiplicand[3];
wire w_pp_11_4 = i_multiplier[11] & i_multiplicand[4];
wire w_pp_11_5 = i_multiplier[11] & i_multiplicand[5];
wire w_pp_11_6 = i_multiplier[11] & i_multiplicand[6];
wire w_pp_11_7 = i_multiplier[11] & i_multiplicand[7];
wire w_pp_11_8 = i_multiplier[11] & i_multiplicand[8];
wire w_pp_11_9 = i_multiplier[11] & i_multiplicand[9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_11_16 = i_multiplier[11] & i_multiplicand[16];
wire w_pp_11_17 = i_multiplier[11] & i_multiplicand[17];
wire w_pp_11_18 = i_multiplier[11] & i_multiplicand[18];
wire w_pp_11_19 = i_multiplier[11] & i_multiplicand[19];
wire w_pp_11_20 = i_multiplier[11] & i_multiplicand[20];
wire w_pp_11_21 = i_multiplier[11] & i_multiplicand[21];
wire w_pp_11_22 = i_multiplier[11] & i_multiplicand[22];
wire w_pp_11_23 = i_multiplier[11] & i_multiplicand[23];
wire w_pp_11_24 = i_multiplier[11] & i_multiplicand[24];
wire w_pp_11_25 = i_multiplier[11] & i_multiplicand[25];
wire w_pp_11_26 = i_multiplier[11] & i_multiplicand[26];
wire w_pp_11_27 = i_multiplier[11] & i_multiplicand[27];
wire w_pp_11_28 = i_multiplier[11] & i_multiplicand[28];
wire w_pp_11_29 = i_multiplier[11] & i_multiplicand[29];
wire w_pp_11_30 = i_multiplier[11] & i_multiplicand[30];
wire w_pp_11_31 = i_multiplier[11] & i_multiplicand[31];
wire w_pp_12_0 = i_multiplier[12] & i_multiplicand[0];
wire w_pp_12_1 = i_multiplier[12] & i_multiplicand[1];
wire w_pp_12_2 = i_multiplier[12] & i_multiplicand[2];
wire w_pp_12_3 = i_multiplier[12] & i_multiplicand[3];
wire w_pp_12_4 = i_multiplier[12] & i_multiplicand[4];
wire w_pp_12_5 = i_multiplier[12] & i_multiplicand[5];
wire w_pp_12_6 = i_multiplier[12] & i_multiplicand[6];
wire w_pp_12_7 = i_multiplier[12] & i_multiplicand[7];
wire w_pp_12_8 = i_multiplier[12] & i_multiplicand[8];
wire w_pp_12_9 = i_multiplier[12] & i_multiplicand[9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_12_16 = i_multiplier[12] & i_multiplicand[16];
wire w_pp_12_17 = i_multiplier[12] & i_multiplicand[17];
wire w_pp_12_18 = i_multiplier[12] & i_multiplicand[18];
wire w_pp_12_19 = i_multiplier[12] & i_multiplicand[19];
wire w_pp_12_20 = i_multiplier[12] & i_multiplicand[20];
wire w_pp_12_21 = i_multiplier[12] & i_multiplicand[21];
wire w_pp_12_22 = i_multiplier[12] & i_multiplicand[22];
wire w_pp_12_23 = i_multiplier[12] & i_multiplicand[23];
wire w_pp_12_24 = i_multiplier[12] & i_multiplicand[24];
wire w_pp_12_25 = i_multiplier[12] & i_multiplicand[25];
wire w_pp_12_26 = i_multiplier[12] & i_multiplicand[26];
wire w_pp_12_27 = i_multiplier[12] & i_multiplicand[27];
wire w_pp_12_28 = i_multiplier[12] & i_multiplicand[28];
wire w_pp_12_29 = i_multiplier[12] & i_multiplicand[29];
wire w_pp_12_30 = i_multiplier[12] & i_multiplicand[30];
wire w_pp_12_31 = i_multiplier[12] & i_multiplicand[31];
wire w_pp_13_0 = i_multiplier[13] & i_multiplicand[0];
wire w_pp_13_1 = i_multiplier[13] & i_multiplicand[1];
wire w_pp_13_2 = i_multiplier[13] & i_multiplicand[2];
wire w_pp_13_3 = i_multiplier[13] & i_multiplicand[3];
wire w_pp_13_4 = i_multiplier[13] & i_multiplicand[4];
wire w_pp_13_5 = i_multiplier[13] & i_multiplicand[5];
wire w_pp_13_6 = i_multiplier[13] & i_multiplicand[6];
wire w_pp_13_7 = i_multiplier[13] & i_multiplicand[7];
wire w_pp_13_8 = i_multiplier[13] & i_multiplicand[8];
wire w_pp_13_9 = i_multiplier[13] & i_multiplicand[9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_13_16 = i_multiplier[13] & i_multiplicand[16];
wire w_pp_13_17 = i_multiplier[13] & i_multiplicand[17];
wire w_pp_13_18 = i_multiplier[13] & i_multiplicand[18];
wire w_pp_13_19 = i_multiplier[13] & i_multiplicand[19];
wire w_pp_13_20 = i_multiplier[13] & i_multiplicand[20];
wire w_pp_13_21 = i_multiplier[13] & i_multiplicand[21];
wire w_pp_13_22 = i_multiplier[13] & i_multiplicand[22];
wire w_pp_13_23 = i_multiplier[13] & i_multiplicand[23];
wire w_pp_13_24 = i_multiplier[13] & i_multiplicand[24];
wire w_pp_13_25 = i_multiplier[13] & i_multiplicand[25];
wire w_pp_13_26 = i_multiplier[13] & i_multiplicand[26];
wire w_pp_13_27 = i_multiplier[13] & i_multiplicand[27];
wire w_pp_13_28 = i_multiplier[13] & i_multiplicand[28];
wire w_pp_13_29 = i_multiplier[13] & i_multiplicand[29];
wire w_pp_13_30 = i_multiplier[13] & i_multiplicand[30];
wire w_pp_13_31 = i_multiplier[13] & i_multiplicand[31];
wire w_pp_14_0 = i_multiplier[14] & i_multiplicand[0];
wire w_pp_14_1 = i_multiplier[14] & i_multiplicand[1];
wire w_pp_14_2 = i_multiplier[14] & i_multiplicand[2];
wire w_pp_14_3 = i_multiplier[14] & i_multiplicand[3];
wire w_pp_14_4 = i_multiplier[14] & i_multiplicand[4];
wire w_pp_14_5 = i_multiplier[14] & i_multiplicand[5];
wire w_pp_14_6 = i_multiplier[14] & i_multiplicand[6];
wire w_pp_14_7 = i_multiplier[14] & i_multiplicand[7];
wire w_pp_14_8 = i_multiplier[14] & i_multiplicand[8];
wire w_pp_14_9 = i_multiplier[14] & i_multiplicand[9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_14_16 = i_multiplier[14] & i_multiplicand[16];
wire w_pp_14_17 = i_multiplier[14] & i_multiplicand[17];
wire w_pp_14_18 = i_multiplier[14] & i_multiplicand[18];
wire w_pp_14_19 = i_multiplier[14] & i_multiplicand[19];
wire w_pp_14_20 = i_multiplier[14] & i_multiplicand[20];
wire w_pp_14_21 = i_multiplier[14] & i_multiplicand[21];
wire w_pp_14_22 = i_multiplier[14] & i_multiplicand[22];
wire w_pp_14_23 = i_multiplier[14] & i_multiplicand[23];
wire w_pp_14_24 = i_multiplier[14] & i_multiplicand[24];
wire w_pp_14_25 = i_multiplier[14] & i_multiplicand[25];
wire w_pp_14_26 = i_multiplier[14] & i_multiplicand[26];
wire w_pp_14_27 = i_multiplier[14] & i_multiplicand[27];
wire w_pp_14_28 = i_multiplier[14] & i_multiplicand[28];
wire w_pp_14_29 = i_multiplier[14] & i_multiplicand[29];
wire w_pp_14_30 = i_multiplier[14] & i_multiplicand[30];
wire w_pp_14_31 = i_multiplier[14] & i_multiplicand[31];
wire w_pp_15_0 = i_multiplier[15] & i_multiplicand[0];
wire w_pp_15_1 = i_multiplier[15] & i_multiplicand[1];
wire w_pp_15_2 = i_multiplier[15] & i_multiplicand[2];
wire w_pp_15_3 = i_multiplier[15] & i_multiplicand[3];
wire w_pp_15_4 = i_multiplier[15] & i_multiplicand[4];
wire w_pp_15_5 = i_multiplier[15] & i_multiplicand[5];
wire w_pp_15_6 = i_multiplier[15] & i_multiplicand[6];
wire w_pp_15_7 = i_multiplier[15] & i_multiplicand[7];
wire w_pp_15_8 = i_multiplier[15] & i_multiplicand[8];
wire w_pp_15_9 = i_multiplier[15] & i_multiplicand[9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];
wire w_pp_15_16 = i_multiplier[15] & i_multiplicand[16];
wire w_pp_15_17 = i_multiplier[15] & i_multiplicand[17];
wire w_pp_15_18 = i_multiplier[15] & i_multiplicand[18];
wire w_pp_15_19 = i_multiplier[15] & i_multiplicand[19];
wire w_pp_15_20 = i_multiplier[15] & i_multiplicand[20];
wire w_pp_15_21 = i_multiplier[15] & i_multiplicand[21];
wire w_pp_15_22 = i_multiplier[15] & i_multiplicand[22];
wire w_pp_15_23 = i_multiplier[15] & i_multiplicand[23];
wire w_pp_15_24 = i_multiplier[15] & i_multiplicand[24];
wire w_pp_15_25 = i_multiplier[15] & i_multiplicand[25];
wire w_pp_15_26 = i_multiplier[15] & i_multiplicand[26];
wire w_pp_15_27 = i_multiplier[15] & i_multiplicand[27];
wire w_pp_15_28 = i_multiplier[15] & i_multiplicand[28];
wire w_pp_15_29 = i_multiplier[15] & i_multiplicand[29];
wire w_pp_15_30 = i_multiplier[15] & i_multiplicand[30];
wire w_pp_15_31 = i_multiplier[15] & i_multiplicand[31];
wire w_pp_16_0 = i_multiplier[16] & i_multiplicand[0];
wire w_pp_16_1 = i_multiplier[16] & i_multiplicand[1];
wire w_pp_16_2 = i_multiplier[16] & i_multiplicand[2];
wire w_pp_16_3 = i_multiplier[16] & i_multiplicand[3];
wire w_pp_16_4 = i_multiplier[16] & i_multiplicand[4];
wire w_pp_16_5 = i_multiplier[16] & i_multiplicand[5];
wire w_pp_16_6 = i_multiplier[16] & i_multiplicand[6];
wire w_pp_16_7 = i_multiplier[16] & i_multiplicand[7];
wire w_pp_16_8 = i_multiplier[16] & i_multiplicand[8];
wire w_pp_16_9 = i_multiplier[16] & i_multiplicand[9];
wire w_pp_16_10 = i_multiplier[16] & i_multiplicand[10];
wire w_pp_16_11 = i_multiplier[16] & i_multiplicand[11];
wire w_pp_16_12 = i_multiplier[16] & i_multiplicand[12];
wire w_pp_16_13 = i_multiplier[16] & i_multiplicand[13];
wire w_pp_16_14 = i_multiplier[16] & i_multiplicand[14];
wire w_pp_16_15 = i_multiplier[16] & i_multiplicand[15];
wire w_pp_16_16 = i_multiplier[16] & i_multiplicand[16];
wire w_pp_16_17 = i_multiplier[16] & i_multiplicand[17];
wire w_pp_16_18 = i_multiplier[16] & i_multiplicand[18];
wire w_pp_16_19 = i_multiplier[16] & i_multiplicand[19];
wire w_pp_16_20 = i_multiplier[16] & i_multiplicand[20];
wire w_pp_16_21 = i_multiplier[16] & i_multiplicand[21];
wire w_pp_16_22 = i_multiplier[16] & i_multiplicand[22];
wire w_pp_16_23 = i_multiplier[16] & i_multiplicand[23];
wire w_pp_16_24 = i_multiplier[16] & i_multiplicand[24];
wire w_pp_16_25 = i_multiplier[16] & i_multiplicand[25];
wire w_pp_16_26 = i_multiplier[16] & i_multiplicand[26];
wire w_pp_16_27 = i_multiplier[16] & i_multiplicand[27];
wire w_pp_16_28 = i_multiplier[16] & i_multiplicand[28];
wire w_pp_16_29 = i_multiplier[16] & i_multiplicand[29];
wire w_pp_16_30 = i_multiplier[16] & i_multiplicand[30];
wire w_pp_16_31 = i_multiplier[16] & i_multiplicand[31];
wire w_pp_17_0 = i_multiplier[17] & i_multiplicand[0];
wire w_pp_17_1 = i_multiplier[17] & i_multiplicand[1];
wire w_pp_17_2 = i_multiplier[17] & i_multiplicand[2];
wire w_pp_17_3 = i_multiplier[17] & i_multiplicand[3];
wire w_pp_17_4 = i_multiplier[17] & i_multiplicand[4];
wire w_pp_17_5 = i_multiplier[17] & i_multiplicand[5];
wire w_pp_17_6 = i_multiplier[17] & i_multiplicand[6];
wire w_pp_17_7 = i_multiplier[17] & i_multiplicand[7];
wire w_pp_17_8 = i_multiplier[17] & i_multiplicand[8];
wire w_pp_17_9 = i_multiplier[17] & i_multiplicand[9];
wire w_pp_17_10 = i_multiplier[17] & i_multiplicand[10];
wire w_pp_17_11 = i_multiplier[17] & i_multiplicand[11];
wire w_pp_17_12 = i_multiplier[17] & i_multiplicand[12];
wire w_pp_17_13 = i_multiplier[17] & i_multiplicand[13];
wire w_pp_17_14 = i_multiplier[17] & i_multiplicand[14];
wire w_pp_17_15 = i_multiplier[17] & i_multiplicand[15];
wire w_pp_17_16 = i_multiplier[17] & i_multiplicand[16];
wire w_pp_17_17 = i_multiplier[17] & i_multiplicand[17];
wire w_pp_17_18 = i_multiplier[17] & i_multiplicand[18];
wire w_pp_17_19 = i_multiplier[17] & i_multiplicand[19];
wire w_pp_17_20 = i_multiplier[17] & i_multiplicand[20];
wire w_pp_17_21 = i_multiplier[17] & i_multiplicand[21];
wire w_pp_17_22 = i_multiplier[17] & i_multiplicand[22];
wire w_pp_17_23 = i_multiplier[17] & i_multiplicand[23];
wire w_pp_17_24 = i_multiplier[17] & i_multiplicand[24];
wire w_pp_17_25 = i_multiplier[17] & i_multiplicand[25];
wire w_pp_17_26 = i_multiplier[17] & i_multiplicand[26];
wire w_pp_17_27 = i_multiplier[17] & i_multiplicand[27];
wire w_pp_17_28 = i_multiplier[17] & i_multiplicand[28];
wire w_pp_17_29 = i_multiplier[17] & i_multiplicand[29];
wire w_pp_17_30 = i_multiplier[17] & i_multiplicand[30];
wire w_pp_17_31 = i_multiplier[17] & i_multiplicand[31];
wire w_pp_18_0 = i_multiplier[18] & i_multiplicand[0];
wire w_pp_18_1 = i_multiplier[18] & i_multiplicand[1];
wire w_pp_18_2 = i_multiplier[18] & i_multiplicand[2];
wire w_pp_18_3 = i_multiplier[18] & i_multiplicand[3];
wire w_pp_18_4 = i_multiplier[18] & i_multiplicand[4];
wire w_pp_18_5 = i_multiplier[18] & i_multiplicand[5];
wire w_pp_18_6 = i_multiplier[18] & i_multiplicand[6];
wire w_pp_18_7 = i_multiplier[18] & i_multiplicand[7];
wire w_pp_18_8 = i_multiplier[18] & i_multiplicand[8];
wire w_pp_18_9 = i_multiplier[18] & i_multiplicand[9];
wire w_pp_18_10 = i_multiplier[18] & i_multiplicand[10];
wire w_pp_18_11 = i_multiplier[18] & i_multiplicand[11];
wire w_pp_18_12 = i_multiplier[18] & i_multiplicand[12];
wire w_pp_18_13 = i_multiplier[18] & i_multiplicand[13];
wire w_pp_18_14 = i_multiplier[18] & i_multiplicand[14];
wire w_pp_18_15 = i_multiplier[18] & i_multiplicand[15];
wire w_pp_18_16 = i_multiplier[18] & i_multiplicand[16];
wire w_pp_18_17 = i_multiplier[18] & i_multiplicand[17];
wire w_pp_18_18 = i_multiplier[18] & i_multiplicand[18];
wire w_pp_18_19 = i_multiplier[18] & i_multiplicand[19];
wire w_pp_18_20 = i_multiplier[18] & i_multiplicand[20];
wire w_pp_18_21 = i_multiplier[18] & i_multiplicand[21];
wire w_pp_18_22 = i_multiplier[18] & i_multiplicand[22];
wire w_pp_18_23 = i_multiplier[18] & i_multiplicand[23];
wire w_pp_18_24 = i_multiplier[18] & i_multiplicand[24];
wire w_pp_18_25 = i_multiplier[18] & i_multiplicand[25];
wire w_pp_18_26 = i_multiplier[18] & i_multiplicand[26];
wire w_pp_18_27 = i_multiplier[18] & i_multiplicand[27];
wire w_pp_18_28 = i_multiplier[18] & i_multiplicand[28];
wire w_pp_18_29 = i_multiplier[18] & i_multiplicand[29];
wire w_pp_18_30 = i_multiplier[18] & i_multiplicand[30];
wire w_pp_18_31 = i_multiplier[18] & i_multiplicand[31];
wire w_pp_19_0 = i_multiplier[19] & i_multiplicand[0];
wire w_pp_19_1 = i_multiplier[19] & i_multiplicand[1];
wire w_pp_19_2 = i_multiplier[19] & i_multiplicand[2];
wire w_pp_19_3 = i_multiplier[19] & i_multiplicand[3];
wire w_pp_19_4 = i_multiplier[19] & i_multiplicand[4];
wire w_pp_19_5 = i_multiplier[19] & i_multiplicand[5];
wire w_pp_19_6 = i_multiplier[19] & i_multiplicand[6];
wire w_pp_19_7 = i_multiplier[19] & i_multiplicand[7];
wire w_pp_19_8 = i_multiplier[19] & i_multiplicand[8];
wire w_pp_19_9 = i_multiplier[19] & i_multiplicand[9];
wire w_pp_19_10 = i_multiplier[19] & i_multiplicand[10];
wire w_pp_19_11 = i_multiplier[19] & i_multiplicand[11];
wire w_pp_19_12 = i_multiplier[19] & i_multiplicand[12];
wire w_pp_19_13 = i_multiplier[19] & i_multiplicand[13];
wire w_pp_19_14 = i_multiplier[19] & i_multiplicand[14];
wire w_pp_19_15 = i_multiplier[19] & i_multiplicand[15];
wire w_pp_19_16 = i_multiplier[19] & i_multiplicand[16];
wire w_pp_19_17 = i_multiplier[19] & i_multiplicand[17];
wire w_pp_19_18 = i_multiplier[19] & i_multiplicand[18];
wire w_pp_19_19 = i_multiplier[19] & i_multiplicand[19];
wire w_pp_19_20 = i_multiplier[19] & i_multiplicand[20];
wire w_pp_19_21 = i_multiplier[19] & i_multiplicand[21];
wire w_pp_19_22 = i_multiplier[19] & i_multiplicand[22];
wire w_pp_19_23 = i_multiplier[19] & i_multiplicand[23];
wire w_pp_19_24 = i_multiplier[19] & i_multiplicand[24];
wire w_pp_19_25 = i_multiplier[19] & i_multiplicand[25];
wire w_pp_19_26 = i_multiplier[19] & i_multiplicand[26];
wire w_pp_19_27 = i_multiplier[19] & i_multiplicand[27];
wire w_pp_19_28 = i_multiplier[19] & i_multiplicand[28];
wire w_pp_19_29 = i_multiplier[19] & i_multiplicand[29];
wire w_pp_19_30 = i_multiplier[19] & i_multiplicand[30];
wire w_pp_19_31 = i_multiplier[19] & i_multiplicand[31];
wire w_pp_20_0 = i_multiplier[20] & i_multiplicand[0];
wire w_pp_20_1 = i_multiplier[20] & i_multiplicand[1];
wire w_pp_20_2 = i_multiplier[20] & i_multiplicand[2];
wire w_pp_20_3 = i_multiplier[20] & i_multiplicand[3];
wire w_pp_20_4 = i_multiplier[20] & i_multiplicand[4];
wire w_pp_20_5 = i_multiplier[20] & i_multiplicand[5];
wire w_pp_20_6 = i_multiplier[20] & i_multiplicand[6];
wire w_pp_20_7 = i_multiplier[20] & i_multiplicand[7];
wire w_pp_20_8 = i_multiplier[20] & i_multiplicand[8];
wire w_pp_20_9 = i_multiplier[20] & i_multiplicand[9];
wire w_pp_20_10 = i_multiplier[20] & i_multiplicand[10];
wire w_pp_20_11 = i_multiplier[20] & i_multiplicand[11];
wire w_pp_20_12 = i_multiplier[20] & i_multiplicand[12];
wire w_pp_20_13 = i_multiplier[20] & i_multiplicand[13];
wire w_pp_20_14 = i_multiplier[20] & i_multiplicand[14];
wire w_pp_20_15 = i_multiplier[20] & i_multiplicand[15];
wire w_pp_20_16 = i_multiplier[20] & i_multiplicand[16];
wire w_pp_20_17 = i_multiplier[20] & i_multiplicand[17];
wire w_pp_20_18 = i_multiplier[20] & i_multiplicand[18];
wire w_pp_20_19 = i_multiplier[20] & i_multiplicand[19];
wire w_pp_20_20 = i_multiplier[20] & i_multiplicand[20];
wire w_pp_20_21 = i_multiplier[20] & i_multiplicand[21];
wire w_pp_20_22 = i_multiplier[20] & i_multiplicand[22];
wire w_pp_20_23 = i_multiplier[20] & i_multiplicand[23];
wire w_pp_20_24 = i_multiplier[20] & i_multiplicand[24];
wire w_pp_20_25 = i_multiplier[20] & i_multiplicand[25];
wire w_pp_20_26 = i_multiplier[20] & i_multiplicand[26];
wire w_pp_20_27 = i_multiplier[20] & i_multiplicand[27];
wire w_pp_20_28 = i_multiplier[20] & i_multiplicand[28];
wire w_pp_20_29 = i_multiplier[20] & i_multiplicand[29];
wire w_pp_20_30 = i_multiplier[20] & i_multiplicand[30];
wire w_pp_20_31 = i_multiplier[20] & i_multiplicand[31];
wire w_pp_21_0 = i_multiplier[21] & i_multiplicand[0];
wire w_pp_21_1 = i_multiplier[21] & i_multiplicand[1];
wire w_pp_21_2 = i_multiplier[21] & i_multiplicand[2];
wire w_pp_21_3 = i_multiplier[21] & i_multiplicand[3];
wire w_pp_21_4 = i_multiplier[21] & i_multiplicand[4];
wire w_pp_21_5 = i_multiplier[21] & i_multiplicand[5];
wire w_pp_21_6 = i_multiplier[21] & i_multiplicand[6];
wire w_pp_21_7 = i_multiplier[21] & i_multiplicand[7];
wire w_pp_21_8 = i_multiplier[21] & i_multiplicand[8];
wire w_pp_21_9 = i_multiplier[21] & i_multiplicand[9];
wire w_pp_21_10 = i_multiplier[21] & i_multiplicand[10];
wire w_pp_21_11 = i_multiplier[21] & i_multiplicand[11];
wire w_pp_21_12 = i_multiplier[21] & i_multiplicand[12];
wire w_pp_21_13 = i_multiplier[21] & i_multiplicand[13];
wire w_pp_21_14 = i_multiplier[21] & i_multiplicand[14];
wire w_pp_21_15 = i_multiplier[21] & i_multiplicand[15];
wire w_pp_21_16 = i_multiplier[21] & i_multiplicand[16];
wire w_pp_21_17 = i_multiplier[21] & i_multiplicand[17];
wire w_pp_21_18 = i_multiplier[21] & i_multiplicand[18];
wire w_pp_21_19 = i_multiplier[21] & i_multiplicand[19];
wire w_pp_21_20 = i_multiplier[21] & i_multiplicand[20];
wire w_pp_21_21 = i_multiplier[21] & i_multiplicand[21];
wire w_pp_21_22 = i_multiplier[21] & i_multiplicand[22];
wire w_pp_21_23 = i_multiplier[21] & i_multiplicand[23];
wire w_pp_21_24 = i_multiplier[21] & i_multiplicand[24];
wire w_pp_21_25 = i_multiplier[21] & i_multiplicand[25];
wire w_pp_21_26 = i_multiplier[21] & i_multiplicand[26];
wire w_pp_21_27 = i_multiplier[21] & i_multiplicand[27];
wire w_pp_21_28 = i_multiplier[21] & i_multiplicand[28];
wire w_pp_21_29 = i_multiplier[21] & i_multiplicand[29];
wire w_pp_21_30 = i_multiplier[21] & i_multiplicand[30];
wire w_pp_21_31 = i_multiplier[21] & i_multiplicand[31];
wire w_pp_22_0 = i_multiplier[22] & i_multiplicand[0];
wire w_pp_22_1 = i_multiplier[22] & i_multiplicand[1];
wire w_pp_22_2 = i_multiplier[22] & i_multiplicand[2];
wire w_pp_22_3 = i_multiplier[22] & i_multiplicand[3];
wire w_pp_22_4 = i_multiplier[22] & i_multiplicand[4];
wire w_pp_22_5 = i_multiplier[22] & i_multiplicand[5];
wire w_pp_22_6 = i_multiplier[22] & i_multiplicand[6];
wire w_pp_22_7 = i_multiplier[22] & i_multiplicand[7];
wire w_pp_22_8 = i_multiplier[22] & i_multiplicand[8];
wire w_pp_22_9 = i_multiplier[22] & i_multiplicand[9];
wire w_pp_22_10 = i_multiplier[22] & i_multiplicand[10];
wire w_pp_22_11 = i_multiplier[22] & i_multiplicand[11];
wire w_pp_22_12 = i_multiplier[22] & i_multiplicand[12];
wire w_pp_22_13 = i_multiplier[22] & i_multiplicand[13];
wire w_pp_22_14 = i_multiplier[22] & i_multiplicand[14];
wire w_pp_22_15 = i_multiplier[22] & i_multiplicand[15];
wire w_pp_22_16 = i_multiplier[22] & i_multiplicand[16];
wire w_pp_22_17 = i_multiplier[22] & i_multiplicand[17];
wire w_pp_22_18 = i_multiplier[22] & i_multiplicand[18];
wire w_pp_22_19 = i_multiplier[22] & i_multiplicand[19];
wire w_pp_22_20 = i_multiplier[22] & i_multiplicand[20];
wire w_pp_22_21 = i_multiplier[22] & i_multiplicand[21];
wire w_pp_22_22 = i_multiplier[22] & i_multiplicand[22];
wire w_pp_22_23 = i_multiplier[22] & i_multiplicand[23];
wire w_pp_22_24 = i_multiplier[22] & i_multiplicand[24];
wire w_pp_22_25 = i_multiplier[22] & i_multiplicand[25];
wire w_pp_22_26 = i_multiplier[22] & i_multiplicand[26];
wire w_pp_22_27 = i_multiplier[22] & i_multiplicand[27];
wire w_pp_22_28 = i_multiplier[22] & i_multiplicand[28];
wire w_pp_22_29 = i_multiplier[22] & i_multiplicand[29];
wire w_pp_22_30 = i_multiplier[22] & i_multiplicand[30];
wire w_pp_22_31 = i_multiplier[22] & i_multiplicand[31];
wire w_pp_23_0 = i_multiplier[23] & i_multiplicand[0];
wire w_pp_23_1 = i_multiplier[23] & i_multiplicand[1];
wire w_pp_23_2 = i_multiplier[23] & i_multiplicand[2];
wire w_pp_23_3 = i_multiplier[23] & i_multiplicand[3];
wire w_pp_23_4 = i_multiplier[23] & i_multiplicand[4];
wire w_pp_23_5 = i_multiplier[23] & i_multiplicand[5];
wire w_pp_23_6 = i_multiplier[23] & i_multiplicand[6];
wire w_pp_23_7 = i_multiplier[23] & i_multiplicand[7];
wire w_pp_23_8 = i_multiplier[23] & i_multiplicand[8];
wire w_pp_23_9 = i_multiplier[23] & i_multiplicand[9];
wire w_pp_23_10 = i_multiplier[23] & i_multiplicand[10];
wire w_pp_23_11 = i_multiplier[23] & i_multiplicand[11];
wire w_pp_23_12 = i_multiplier[23] & i_multiplicand[12];
wire w_pp_23_13 = i_multiplier[23] & i_multiplicand[13];
wire w_pp_23_14 = i_multiplier[23] & i_multiplicand[14];
wire w_pp_23_15 = i_multiplier[23] & i_multiplicand[15];
wire w_pp_23_16 = i_multiplier[23] & i_multiplicand[16];
wire w_pp_23_17 = i_multiplier[23] & i_multiplicand[17];
wire w_pp_23_18 = i_multiplier[23] & i_multiplicand[18];
wire w_pp_23_19 = i_multiplier[23] & i_multiplicand[19];
wire w_pp_23_20 = i_multiplier[23] & i_multiplicand[20];
wire w_pp_23_21 = i_multiplier[23] & i_multiplicand[21];
wire w_pp_23_22 = i_multiplier[23] & i_multiplicand[22];
wire w_pp_23_23 = i_multiplier[23] & i_multiplicand[23];
wire w_pp_23_24 = i_multiplier[23] & i_multiplicand[24];
wire w_pp_23_25 = i_multiplier[23] & i_multiplicand[25];
wire w_pp_23_26 = i_multiplier[23] & i_multiplicand[26];
wire w_pp_23_27 = i_multiplier[23] & i_multiplicand[27];
wire w_pp_23_28 = i_multiplier[23] & i_multiplicand[28];
wire w_pp_23_29 = i_multiplier[23] & i_multiplicand[29];
wire w_pp_23_30 = i_multiplier[23] & i_multiplicand[30];
wire w_pp_23_31 = i_multiplier[23] & i_multiplicand[31];
wire w_pp_24_0 = i_multiplier[24] & i_multiplicand[0];
wire w_pp_24_1 = i_multiplier[24] & i_multiplicand[1];
wire w_pp_24_2 = i_multiplier[24] & i_multiplicand[2];
wire w_pp_24_3 = i_multiplier[24] & i_multiplicand[3];
wire w_pp_24_4 = i_multiplier[24] & i_multiplicand[4];
wire w_pp_24_5 = i_multiplier[24] & i_multiplicand[5];
wire w_pp_24_6 = i_multiplier[24] & i_multiplicand[6];
wire w_pp_24_7 = i_multiplier[24] & i_multiplicand[7];
wire w_pp_24_8 = i_multiplier[24] & i_multiplicand[8];
wire w_pp_24_9 = i_multiplier[24] & i_multiplicand[9];
wire w_pp_24_10 = i_multiplier[24] & i_multiplicand[10];
wire w_pp_24_11 = i_multiplier[24] & i_multiplicand[11];
wire w_pp_24_12 = i_multiplier[24] & i_multiplicand[12];
wire w_pp_24_13 = i_multiplier[24] & i_multiplicand[13];
wire w_pp_24_14 = i_multiplier[24] & i_multiplicand[14];
wire w_pp_24_15 = i_multiplier[24] & i_multiplicand[15];
wire w_pp_24_16 = i_multiplier[24] & i_multiplicand[16];
wire w_pp_24_17 = i_multiplier[24] & i_multiplicand[17];
wire w_pp_24_18 = i_multiplier[24] & i_multiplicand[18];
wire w_pp_24_19 = i_multiplier[24] & i_multiplicand[19];
wire w_pp_24_20 = i_multiplier[24] & i_multiplicand[20];
wire w_pp_24_21 = i_multiplier[24] & i_multiplicand[21];
wire w_pp_24_22 = i_multiplier[24] & i_multiplicand[22];
wire w_pp_24_23 = i_multiplier[24] & i_multiplicand[23];
wire w_pp_24_24 = i_multiplier[24] & i_multiplicand[24];
wire w_pp_24_25 = i_multiplier[24] & i_multiplicand[25];
wire w_pp_24_26 = i_multiplier[24] & i_multiplicand[26];
wire w_pp_24_27 = i_multiplier[24] & i_multiplicand[27];
wire w_pp_24_28 = i_multiplier[24] & i_multiplicand[28];
wire w_pp_24_29 = i_multiplier[24] & i_multiplicand[29];
wire w_pp_24_30 = i_multiplier[24] & i_multiplicand[30];
wire w_pp_24_31 = i_multiplier[24] & i_multiplicand[31];
wire w_pp_25_0 = i_multiplier[25] & i_multiplicand[0];
wire w_pp_25_1 = i_multiplier[25] & i_multiplicand[1];
wire w_pp_25_2 = i_multiplier[25] & i_multiplicand[2];
wire w_pp_25_3 = i_multiplier[25] & i_multiplicand[3];
wire w_pp_25_4 = i_multiplier[25] & i_multiplicand[4];
wire w_pp_25_5 = i_multiplier[25] & i_multiplicand[5];
wire w_pp_25_6 = i_multiplier[25] & i_multiplicand[6];
wire w_pp_25_7 = i_multiplier[25] & i_multiplicand[7];
wire w_pp_25_8 = i_multiplier[25] & i_multiplicand[8];
wire w_pp_25_9 = i_multiplier[25] & i_multiplicand[9];
wire w_pp_25_10 = i_multiplier[25] & i_multiplicand[10];
wire w_pp_25_11 = i_multiplier[25] & i_multiplicand[11];
wire w_pp_25_12 = i_multiplier[25] & i_multiplicand[12];
wire w_pp_25_13 = i_multiplier[25] & i_multiplicand[13];
wire w_pp_25_14 = i_multiplier[25] & i_multiplicand[14];
wire w_pp_25_15 = i_multiplier[25] & i_multiplicand[15];
wire w_pp_25_16 = i_multiplier[25] & i_multiplicand[16];
wire w_pp_25_17 = i_multiplier[25] & i_multiplicand[17];
wire w_pp_25_18 = i_multiplier[25] & i_multiplicand[18];
wire w_pp_25_19 = i_multiplier[25] & i_multiplicand[19];
wire w_pp_25_20 = i_multiplier[25] & i_multiplicand[20];
wire w_pp_25_21 = i_multiplier[25] & i_multiplicand[21];
wire w_pp_25_22 = i_multiplier[25] & i_multiplicand[22];
wire w_pp_25_23 = i_multiplier[25] & i_multiplicand[23];
wire w_pp_25_24 = i_multiplier[25] & i_multiplicand[24];
wire w_pp_25_25 = i_multiplier[25] & i_multiplicand[25];
wire w_pp_25_26 = i_multiplier[25] & i_multiplicand[26];
wire w_pp_25_27 = i_multiplier[25] & i_multiplicand[27];
wire w_pp_25_28 = i_multiplier[25] & i_multiplicand[28];
wire w_pp_25_29 = i_multiplier[25] & i_multiplicand[29];
wire w_pp_25_30 = i_multiplier[25] & i_multiplicand[30];
wire w_pp_25_31 = i_multiplier[25] & i_multiplicand[31];
wire w_pp_26_0 = i_multiplier[26] & i_multiplicand[0];
wire w_pp_26_1 = i_multiplier[26] & i_multiplicand[1];
wire w_pp_26_2 = i_multiplier[26] & i_multiplicand[2];
wire w_pp_26_3 = i_multiplier[26] & i_multiplicand[3];
wire w_pp_26_4 = i_multiplier[26] & i_multiplicand[4];
wire w_pp_26_5 = i_multiplier[26] & i_multiplicand[5];
wire w_pp_26_6 = i_multiplier[26] & i_multiplicand[6];
wire w_pp_26_7 = i_multiplier[26] & i_multiplicand[7];
wire w_pp_26_8 = i_multiplier[26] & i_multiplicand[8];
wire w_pp_26_9 = i_multiplier[26] & i_multiplicand[9];
wire w_pp_26_10 = i_multiplier[26] & i_multiplicand[10];
wire w_pp_26_11 = i_multiplier[26] & i_multiplicand[11];
wire w_pp_26_12 = i_multiplier[26] & i_multiplicand[12];
wire w_pp_26_13 = i_multiplier[26] & i_multiplicand[13];
wire w_pp_26_14 = i_multiplier[26] & i_multiplicand[14];
wire w_pp_26_15 = i_multiplier[26] & i_multiplicand[15];
wire w_pp_26_16 = i_multiplier[26] & i_multiplicand[16];
wire w_pp_26_17 = i_multiplier[26] & i_multiplicand[17];
wire w_pp_26_18 = i_multiplier[26] & i_multiplicand[18];
wire w_pp_26_19 = i_multiplier[26] & i_multiplicand[19];
wire w_pp_26_20 = i_multiplier[26] & i_multiplicand[20];
wire w_pp_26_21 = i_multiplier[26] & i_multiplicand[21];
wire w_pp_26_22 = i_multiplier[26] & i_multiplicand[22];
wire w_pp_26_23 = i_multiplier[26] & i_multiplicand[23];
wire w_pp_26_24 = i_multiplier[26] & i_multiplicand[24];
wire w_pp_26_25 = i_multiplier[26] & i_multiplicand[25];
wire w_pp_26_26 = i_multiplier[26] & i_multiplicand[26];
wire w_pp_26_27 = i_multiplier[26] & i_multiplicand[27];
wire w_pp_26_28 = i_multiplier[26] & i_multiplicand[28];
wire w_pp_26_29 = i_multiplier[26] & i_multiplicand[29];
wire w_pp_26_30 = i_multiplier[26] & i_multiplicand[30];
wire w_pp_26_31 = i_multiplier[26] & i_multiplicand[31];
wire w_pp_27_0 = i_multiplier[27] & i_multiplicand[0];
wire w_pp_27_1 = i_multiplier[27] & i_multiplicand[1];
wire w_pp_27_2 = i_multiplier[27] & i_multiplicand[2];
wire w_pp_27_3 = i_multiplier[27] & i_multiplicand[3];
wire w_pp_27_4 = i_multiplier[27] & i_multiplicand[4];
wire w_pp_27_5 = i_multiplier[27] & i_multiplicand[5];
wire w_pp_27_6 = i_multiplier[27] & i_multiplicand[6];
wire w_pp_27_7 = i_multiplier[27] & i_multiplicand[7];
wire w_pp_27_8 = i_multiplier[27] & i_multiplicand[8];
wire w_pp_27_9 = i_multiplier[27] & i_multiplicand[9];
wire w_pp_27_10 = i_multiplier[27] & i_multiplicand[10];
wire w_pp_27_11 = i_multiplier[27] & i_multiplicand[11];
wire w_pp_27_12 = i_multiplier[27] & i_multiplicand[12];
wire w_pp_27_13 = i_multiplier[27] & i_multiplicand[13];
wire w_pp_27_14 = i_multiplier[27] & i_multiplicand[14];
wire w_pp_27_15 = i_multiplier[27] & i_multiplicand[15];
wire w_pp_27_16 = i_multiplier[27] & i_multiplicand[16];
wire w_pp_27_17 = i_multiplier[27] & i_multiplicand[17];
wire w_pp_27_18 = i_multiplier[27] & i_multiplicand[18];
wire w_pp_27_19 = i_multiplier[27] & i_multiplicand[19];
wire w_pp_27_20 = i_multiplier[27] & i_multiplicand[20];
wire w_pp_27_21 = i_multiplier[27] & i_multiplicand[21];
wire w_pp_27_22 = i_multiplier[27] & i_multiplicand[22];
wire w_pp_27_23 = i_multiplier[27] & i_multiplicand[23];
wire w_pp_27_24 = i_multiplier[27] & i_multiplicand[24];
wire w_pp_27_25 = i_multiplier[27] & i_multiplicand[25];
wire w_pp_27_26 = i_multiplier[27] & i_multiplicand[26];
wire w_pp_27_27 = i_multiplier[27] & i_multiplicand[27];
wire w_pp_27_28 = i_multiplier[27] & i_multiplicand[28];
wire w_pp_27_29 = i_multiplier[27] & i_multiplicand[29];
wire w_pp_27_30 = i_multiplier[27] & i_multiplicand[30];
wire w_pp_27_31 = i_multiplier[27] & i_multiplicand[31];
wire w_pp_28_0 = i_multiplier[28] & i_multiplicand[0];
wire w_pp_28_1 = i_multiplier[28] & i_multiplicand[1];
wire w_pp_28_2 = i_multiplier[28] & i_multiplicand[2];
wire w_pp_28_3 = i_multiplier[28] & i_multiplicand[3];
wire w_pp_28_4 = i_multiplier[28] & i_multiplicand[4];
wire w_pp_28_5 = i_multiplier[28] & i_multiplicand[5];
wire w_pp_28_6 = i_multiplier[28] & i_multiplicand[6];
wire w_pp_28_7 = i_multiplier[28] & i_multiplicand[7];
wire w_pp_28_8 = i_multiplier[28] & i_multiplicand[8];
wire w_pp_28_9 = i_multiplier[28] & i_multiplicand[9];
wire w_pp_28_10 = i_multiplier[28] & i_multiplicand[10];
wire w_pp_28_11 = i_multiplier[28] & i_multiplicand[11];
wire w_pp_28_12 = i_multiplier[28] & i_multiplicand[12];
wire w_pp_28_13 = i_multiplier[28] & i_multiplicand[13];
wire w_pp_28_14 = i_multiplier[28] & i_multiplicand[14];
wire w_pp_28_15 = i_multiplier[28] & i_multiplicand[15];
wire w_pp_28_16 = i_multiplier[28] & i_multiplicand[16];
wire w_pp_28_17 = i_multiplier[28] & i_multiplicand[17];
wire w_pp_28_18 = i_multiplier[28] & i_multiplicand[18];
wire w_pp_28_19 = i_multiplier[28] & i_multiplicand[19];
wire w_pp_28_20 = i_multiplier[28] & i_multiplicand[20];
wire w_pp_28_21 = i_multiplier[28] & i_multiplicand[21];
wire w_pp_28_22 = i_multiplier[28] & i_multiplicand[22];
wire w_pp_28_23 = i_multiplier[28] & i_multiplicand[23];
wire w_pp_28_24 = i_multiplier[28] & i_multiplicand[24];
wire w_pp_28_25 = i_multiplier[28] & i_multiplicand[25];
wire w_pp_28_26 = i_multiplier[28] & i_multiplicand[26];
wire w_pp_28_27 = i_multiplier[28] & i_multiplicand[27];
wire w_pp_28_28 = i_multiplier[28] & i_multiplicand[28];
wire w_pp_28_29 = i_multiplier[28] & i_multiplicand[29];
wire w_pp_28_30 = i_multiplier[28] & i_multiplicand[30];
wire w_pp_28_31 = i_multiplier[28] & i_multiplicand[31];
wire w_pp_29_0 = i_multiplier[29] & i_multiplicand[0];
wire w_pp_29_1 = i_multiplier[29] & i_multiplicand[1];
wire w_pp_29_2 = i_multiplier[29] & i_multiplicand[2];
wire w_pp_29_3 = i_multiplier[29] & i_multiplicand[3];
wire w_pp_29_4 = i_multiplier[29] & i_multiplicand[4];
wire w_pp_29_5 = i_multiplier[29] & i_multiplicand[5];
wire w_pp_29_6 = i_multiplier[29] & i_multiplicand[6];
wire w_pp_29_7 = i_multiplier[29] & i_multiplicand[7];
wire w_pp_29_8 = i_multiplier[29] & i_multiplicand[8];
wire w_pp_29_9 = i_multiplier[29] & i_multiplicand[9];
wire w_pp_29_10 = i_multiplier[29] & i_multiplicand[10];
wire w_pp_29_11 = i_multiplier[29] & i_multiplicand[11];
wire w_pp_29_12 = i_multiplier[29] & i_multiplicand[12];
wire w_pp_29_13 = i_multiplier[29] & i_multiplicand[13];
wire w_pp_29_14 = i_multiplier[29] & i_multiplicand[14];
wire w_pp_29_15 = i_multiplier[29] & i_multiplicand[15];
wire w_pp_29_16 = i_multiplier[29] & i_multiplicand[16];
wire w_pp_29_17 = i_multiplier[29] & i_multiplicand[17];
wire w_pp_29_18 = i_multiplier[29] & i_multiplicand[18];
wire w_pp_29_19 = i_multiplier[29] & i_multiplicand[19];
wire w_pp_29_20 = i_multiplier[29] & i_multiplicand[20];
wire w_pp_29_21 = i_multiplier[29] & i_multiplicand[21];
wire w_pp_29_22 = i_multiplier[29] & i_multiplicand[22];
wire w_pp_29_23 = i_multiplier[29] & i_multiplicand[23];
wire w_pp_29_24 = i_multiplier[29] & i_multiplicand[24];
wire w_pp_29_25 = i_multiplier[29] & i_multiplicand[25];
wire w_pp_29_26 = i_multiplier[29] & i_multiplicand[26];
wire w_pp_29_27 = i_multiplier[29] & i_multiplicand[27];
wire w_pp_29_28 = i_multiplier[29] & i_multiplicand[28];
wire w_pp_29_29 = i_multiplier[29] & i_multiplicand[29];
wire w_pp_29_30 = i_multiplier[29] & i_multiplicand[30];
wire w_pp_29_31 = i_multiplier[29] & i_multiplicand[31];
wire w_pp_30_0 = i_multiplier[30] & i_multiplicand[0];
wire w_pp_30_1 = i_multiplier[30] & i_multiplicand[1];
wire w_pp_30_2 = i_multiplier[30] & i_multiplicand[2];
wire w_pp_30_3 = i_multiplier[30] & i_multiplicand[3];
wire w_pp_30_4 = i_multiplier[30] & i_multiplicand[4];
wire w_pp_30_5 = i_multiplier[30] & i_multiplicand[5];
wire w_pp_30_6 = i_multiplier[30] & i_multiplicand[6];
wire w_pp_30_7 = i_multiplier[30] & i_multiplicand[7];
wire w_pp_30_8 = i_multiplier[30] & i_multiplicand[8];
wire w_pp_30_9 = i_multiplier[30] & i_multiplicand[9];
wire w_pp_30_10 = i_multiplier[30] & i_multiplicand[10];
wire w_pp_30_11 = i_multiplier[30] & i_multiplicand[11];
wire w_pp_30_12 = i_multiplier[30] & i_multiplicand[12];
wire w_pp_30_13 = i_multiplier[30] & i_multiplicand[13];
wire w_pp_30_14 = i_multiplier[30] & i_multiplicand[14];
wire w_pp_30_15 = i_multiplier[30] & i_multiplicand[15];
wire w_pp_30_16 = i_multiplier[30] & i_multiplicand[16];
wire w_pp_30_17 = i_multiplier[30] & i_multiplicand[17];
wire w_pp_30_18 = i_multiplier[30] & i_multiplicand[18];
wire w_pp_30_19 = i_multiplier[30] & i_multiplicand[19];
wire w_pp_30_20 = i_multiplier[30] & i_multiplicand[20];
wire w_pp_30_21 = i_multiplier[30] & i_multiplicand[21];
wire w_pp_30_22 = i_multiplier[30] & i_multiplicand[22];
wire w_pp_30_23 = i_multiplier[30] & i_multiplicand[23];
wire w_pp_30_24 = i_multiplier[30] & i_multiplicand[24];
wire w_pp_30_25 = i_multiplier[30] & i_multiplicand[25];
wire w_pp_30_26 = i_multiplier[30] & i_multiplicand[26];
wire w_pp_30_27 = i_multiplier[30] & i_multiplicand[27];
wire w_pp_30_28 = i_multiplier[30] & i_multiplicand[28];
wire w_pp_30_29 = i_multiplier[30] & i_multiplicand[29];
wire w_pp_30_30 = i_multiplier[30] & i_multiplicand[30];
wire w_pp_30_31 = i_multiplier[30] & i_multiplicand[31];
wire w_pp_31_0 = i_multiplier[31] & i_multiplicand[0];
wire w_pp_31_1 = i_multiplier[31] & i_multiplicand[1];
wire w_pp_31_2 = i_multiplier[31] & i_multiplicand[2];
wire w_pp_31_3 = i_multiplier[31] & i_multiplicand[3];
wire w_pp_31_4 = i_multiplier[31] & i_multiplicand[4];
wire w_pp_31_5 = i_multiplier[31] & i_multiplicand[5];
wire w_pp_31_6 = i_multiplier[31] & i_multiplicand[6];
wire w_pp_31_7 = i_multiplier[31] & i_multiplicand[7];
wire w_pp_31_8 = i_multiplier[31] & i_multiplicand[8];
wire w_pp_31_9 = i_multiplier[31] & i_multiplicand[9];
wire w_pp_31_10 = i_multiplier[31] & i_multiplicand[10];
wire w_pp_31_11 = i_multiplier[31] & i_multiplicand[11];
wire w_pp_31_12 = i_multiplier[31] & i_multiplicand[12];
wire w_pp_31_13 = i_multiplier[31] & i_multiplicand[13];
wire w_pp_31_14 = i_multiplier[31] & i_multiplicand[14];
wire w_pp_31_15 = i_multiplier[31] & i_multiplicand[15];
wire w_pp_31_16 = i_multiplier[31] & i_multiplicand[16];
wire w_pp_31_17 = i_multiplier[31] & i_multiplicand[17];
wire w_pp_31_18 = i_multiplier[31] & i_multiplicand[18];
wire w_pp_31_19 = i_multiplier[31] & i_multiplicand[19];
wire w_pp_31_20 = i_multiplier[31] & i_multiplicand[20];
wire w_pp_31_21 = i_multiplier[31] & i_multiplicand[21];
wire w_pp_31_22 = i_multiplier[31] & i_multiplicand[22];
wire w_pp_31_23 = i_multiplier[31] & i_multiplicand[23];
wire w_pp_31_24 = i_multiplier[31] & i_multiplicand[24];
wire w_pp_31_25 = i_multiplier[31] & i_multiplicand[25];
wire w_pp_31_26 = i_multiplier[31] & i_multiplicand[26];
wire w_pp_31_27 = i_multiplier[31] & i_multiplicand[27];
wire w_pp_31_28 = i_multiplier[31] & i_multiplicand[28];
wire w_pp_31_29 = i_multiplier[31] & i_multiplicand[29];
wire w_pp_31_30 = i_multiplier[31] & i_multiplicand[30];
wire w_pp_31_31 = i_multiplier[31] & i_multiplicand[31];

// Partial products reduction using Wallace tree
wire w_sum_1_2, w_carry_1_2;
math_adder_half HA_1_2(.i_a(w_pp_0_1), .i_b(w_pp_1_0), .ow_sum(w_sum_1_2), .ow_c(w_carry_1_2));
wire w_sum_2_4, w_carry_2_4;
math_adder_carry_save CSA_2_4(.i_a(w_pp_0_2), .i_b(w_pp_1_1), .i_c(w_pp_2_0), .ow_sum(w_sum_2_4), .ow_c(w_carry_2_4));
wire w_sum_2_2, w_carry_2_2;
math_adder_half HA_2_2(.i_a(w_carry_1_2), .i_b(w_sum_2_4), .ow_sum(w_sum_2_2), .ow_c(w_carry_2_2));
wire w_sum_3_6, w_carry_3_6;
math_adder_carry_save CSA_3_6(.i_a(w_pp_0_3), .i_b(w_pp_1_2), .i_c(w_pp_2_1), .ow_sum(w_sum_3_6), .ow_c(w_carry_3_6));
wire w_sum_3_4, w_carry_3_4;
math_adder_carry_save CSA_3_4(.i_a(w_pp_3_0), .i_b(w_carry_2_4), .i_c(w_carry_2_2), .ow_sum(w_sum_3_4), .ow_c(w_carry_3_4));
wire w_sum_3_2, w_carry_3_2;
math_adder_half HA_3_2(.i_a(w_sum_3_6), .i_b(w_sum_3_4), .ow_sum(w_sum_3_2), .ow_c(w_carry_3_2));
wire w_sum_4_8, w_carry_4_8;
math_adder_carry_save CSA_4_8(.i_a(w_pp_0_4), .i_b(w_pp_1_3), .i_c(w_pp_2_2), .ow_sum(w_sum_4_8), .ow_c(w_carry_4_8));
wire w_sum_4_6, w_carry_4_6;
math_adder_carry_save CSA_4_6(.i_a(w_pp_3_1), .i_b(w_pp_4_0), .i_c(w_carry_3_6), .ow_sum(w_sum_4_6), .ow_c(w_carry_4_6));
wire w_sum_4_4, w_carry_4_4;
math_adder_carry_save CSA_4_4(.i_a(w_carry_3_4), .i_b(w_carry_3_2), .i_c(w_sum_4_8), .ow_sum(w_sum_4_4), .ow_c(w_carry_4_4));
wire w_sum_4_2, w_carry_4_2;
math_adder_half HA_4_2(.i_a(w_sum_4_6), .i_b(w_sum_4_4), .ow_sum(w_sum_4_2), .ow_c(w_carry_4_2));
wire w_sum_5_10, w_carry_5_10;
math_adder_carry_save CSA_5_10(.i_a(w_pp_0_5), .i_b(w_pp_1_4), .i_c(w_pp_2_3), .ow_sum(w_sum_5_10), .ow_c(w_carry_5_10));
wire w_sum_5_8, w_carry_5_8;
math_adder_carry_save CSA_5_8(.i_a(w_pp_3_2), .i_b(w_pp_4_1), .i_c(w_pp_5_0), .ow_sum(w_sum_5_8), .ow_c(w_carry_5_8));
wire w_sum_5_6, w_carry_5_6;
math_adder_carry_save CSA_5_6(.i_a(w_carry_4_8), .i_b(w_carry_4_6), .i_c(w_carry_4_4), .ow_sum(w_sum_5_6), .ow_c(w_carry_5_6));
wire w_sum_5_4, w_carry_5_4;
math_adder_carry_save CSA_5_4(.i_a(w_carry_4_2), .i_b(w_sum_5_10), .i_c(w_sum_5_8), .ow_sum(w_sum_5_4), .ow_c(w_carry_5_4));
wire w_sum_5_2, w_carry_5_2;
math_adder_half HA_5_2(.i_a(w_sum_5_6), .i_b(w_sum_5_4), .ow_sum(w_sum_5_2), .ow_c(w_carry_5_2));
wire w_sum_6_12, w_carry_6_12;
math_adder_carry_save CSA_6_12(.i_a(w_pp_0_6), .i_b(w_pp_1_5), .i_c(w_pp_2_4), .ow_sum(w_sum_6_12), .ow_c(w_carry_6_12));
wire w_sum_6_10, w_carry_6_10;
math_adder_carry_save CSA_6_10(.i_a(w_pp_3_3), .i_b(w_pp_4_2), .i_c(w_pp_5_1), .ow_sum(w_sum_6_10), .ow_c(w_carry_6_10));
wire w_sum_6_8, w_carry_6_8;
math_adder_carry_save CSA_6_8(.i_a(w_pp_6_0), .i_b(w_carry_5_10), .i_c(w_carry_5_8), .ow_sum(w_sum_6_8), .ow_c(w_carry_6_8));
wire w_sum_6_6, w_carry_6_6;
math_adder_carry_save CSA_6_6(.i_a(w_carry_5_6), .i_b(w_carry_5_4), .i_c(w_carry_5_2), .ow_sum(w_sum_6_6), .ow_c(w_carry_6_6));
wire w_sum_6_4, w_carry_6_4;
math_adder_carry_save CSA_6_4(.i_a(w_sum_6_12), .i_b(w_sum_6_10), .i_c(w_sum_6_8), .ow_sum(w_sum_6_4), .ow_c(w_carry_6_4));
wire w_sum_6_2, w_carry_6_2;
math_adder_half HA_6_2(.i_a(w_sum_6_6), .i_b(w_sum_6_4), .ow_sum(w_sum_6_2), .ow_c(w_carry_6_2));
wire w_sum_7_14, w_carry_7_14;
math_adder_carry_save CSA_7_14(.i_a(w_pp_0_7), .i_b(w_pp_1_6), .i_c(w_pp_2_5), .ow_sum(w_sum_7_14), .ow_c(w_carry_7_14));
wire w_sum_7_12, w_carry_7_12;
math_adder_carry_save CSA_7_12(.i_a(w_pp_3_4), .i_b(w_pp_4_3), .i_c(w_pp_5_2), .ow_sum(w_sum_7_12), .ow_c(w_carry_7_12));
wire w_sum_7_10, w_carry_7_10;
math_adder_carry_save CSA_7_10(.i_a(w_pp_6_1), .i_b(w_pp_7_0), .i_c(w_carry_6_12), .ow_sum(w_sum_7_10), .ow_c(w_carry_7_10));
wire w_sum_7_8, w_carry_7_8;
math_adder_carry_save CSA_7_8(.i_a(w_carry_6_10), .i_b(w_carry_6_8), .i_c(w_carry_6_6), .ow_sum(w_sum_7_8), .ow_c(w_carry_7_8));
wire w_sum_7_6, w_carry_7_6;
math_adder_carry_save CSA_7_6(.i_a(w_carry_6_4), .i_b(w_carry_6_2), .i_c(w_sum_7_14), .ow_sum(w_sum_7_6), .ow_c(w_carry_7_6));
wire w_sum_7_4, w_carry_7_4;
math_adder_carry_save CSA_7_4(.i_a(w_sum_7_12), .i_b(w_sum_7_10), .i_c(w_sum_7_8), .ow_sum(w_sum_7_4), .ow_c(w_carry_7_4));
wire w_sum_7_2, w_carry_7_2;
math_adder_half HA_7_2(.i_a(w_sum_7_6), .i_b(w_sum_7_4), .ow_sum(w_sum_7_2), .ow_c(w_carry_7_2));
wire w_sum_8_16, w_carry_8_16;
math_adder_carry_save CSA_8_16(.i_a(w_pp_0_8), .i_b(w_pp_1_7), .i_c(w_pp_2_6), .ow_sum(w_sum_8_16), .ow_c(w_carry_8_16));
wire w_sum_8_14, w_carry_8_14;
math_adder_carry_save CSA_8_14(.i_a(w_pp_3_5), .i_b(w_pp_4_4), .i_c(w_pp_5_3), .ow_sum(w_sum_8_14), .ow_c(w_carry_8_14));
wire w_sum_8_12, w_carry_8_12;
math_adder_carry_save CSA_8_12(.i_a(w_pp_6_2), .i_b(w_pp_7_1), .i_c(w_pp_8_0), .ow_sum(w_sum_8_12), .ow_c(w_carry_8_12));
wire w_sum_8_10, w_carry_8_10;
math_adder_carry_save CSA_8_10(.i_a(w_carry_7_14), .i_b(w_carry_7_12), .i_c(w_carry_7_10), .ow_sum(w_sum_8_10), .ow_c(w_carry_8_10));
wire w_sum_8_8, w_carry_8_8;
math_adder_carry_save CSA_8_8(.i_a(w_carry_7_8), .i_b(w_carry_7_6), .i_c(w_carry_7_4), .ow_sum(w_sum_8_8), .ow_c(w_carry_8_8));
wire w_sum_8_6, w_carry_8_6;
math_adder_carry_save CSA_8_6(.i_a(w_carry_7_2), .i_b(w_sum_8_16), .i_c(w_sum_8_14), .ow_sum(w_sum_8_6), .ow_c(w_carry_8_6));
wire w_sum_8_4, w_carry_8_4;
math_adder_carry_save CSA_8_4(.i_a(w_sum_8_12), .i_b(w_sum_8_10), .i_c(w_sum_8_8), .ow_sum(w_sum_8_4), .ow_c(w_carry_8_4));
wire w_sum_8_2, w_carry_8_2;
math_adder_half HA_8_2(.i_a(w_sum_8_6), .i_b(w_sum_8_4), .ow_sum(w_sum_8_2), .ow_c(w_carry_8_2));
wire w_sum_9_18, w_carry_9_18;
math_adder_carry_save CSA_9_18(.i_a(w_pp_0_9), .i_b(w_pp_1_8), .i_c(w_pp_2_7), .ow_sum(w_sum_9_18), .ow_c(w_carry_9_18));
wire w_sum_9_16, w_carry_9_16;
math_adder_carry_save CSA_9_16(.i_a(w_pp_3_6), .i_b(w_pp_4_5), .i_c(w_pp_5_4), .ow_sum(w_sum_9_16), .ow_c(w_carry_9_16));
wire w_sum_9_14, w_carry_9_14;
math_adder_carry_save CSA_9_14(.i_a(w_pp_6_3), .i_b(w_pp_7_2), .i_c(w_pp_8_1), .ow_sum(w_sum_9_14), .ow_c(w_carry_9_14));
wire w_sum_9_12, w_carry_9_12;
math_adder_carry_save CSA_9_12(.i_a(w_pp_9_0), .i_b(w_carry_8_16), .i_c(w_carry_8_14), .ow_sum(w_sum_9_12), .ow_c(w_carry_9_12));
wire w_sum_9_10, w_carry_9_10;
math_adder_carry_save CSA_9_10(.i_a(w_carry_8_12), .i_b(w_carry_8_10), .i_c(w_carry_8_8), .ow_sum(w_sum_9_10), .ow_c(w_carry_9_10));
wire w_sum_9_8, w_carry_9_8;
math_adder_carry_save CSA_9_8(.i_a(w_carry_8_6), .i_b(w_carry_8_4), .i_c(w_carry_8_2), .ow_sum(w_sum_9_8), .ow_c(w_carry_9_8));
wire w_sum_9_6, w_carry_9_6;
math_adder_carry_save CSA_9_6(.i_a(w_sum_9_18), .i_b(w_sum_9_16), .i_c(w_sum_9_14), .ow_sum(w_sum_9_6), .ow_c(w_carry_9_6));
wire w_sum_9_4, w_carry_9_4;
math_adder_carry_save CSA_9_4(.i_a(w_sum_9_12), .i_b(w_sum_9_10), .i_c(w_sum_9_8), .ow_sum(w_sum_9_4), .ow_c(w_carry_9_4));
wire w_sum_9_2, w_carry_9_2;
math_adder_half HA_9_2(.i_a(w_sum_9_6), .i_b(w_sum_9_4), .ow_sum(w_sum_9_2), .ow_c(w_carry_9_2));
wire w_sum_10_20, w_carry_10_20;
math_adder_carry_save CSA_10_20(.i_a(w_pp_0_10), .i_b(w_pp_1_9), .i_c(w_pp_2_8), .ow_sum(w_sum_10_20), .ow_c(w_carry_10_20));
wire w_sum_10_18, w_carry_10_18;
math_adder_carry_save CSA_10_18(.i_a(w_pp_3_7), .i_b(w_pp_4_6), .i_c(w_pp_5_5), .ow_sum(w_sum_10_18), .ow_c(w_carry_10_18));
wire w_sum_10_16, w_carry_10_16;
math_adder_carry_save CSA_10_16(.i_a(w_pp_6_4), .i_b(w_pp_7_3), .i_c(w_pp_8_2), .ow_sum(w_sum_10_16), .ow_c(w_carry_10_16));
wire w_sum_10_14, w_carry_10_14;
math_adder_carry_save CSA_10_14(.i_a(w_pp_9_1), .i_b(w_pp_10_0), .i_c(w_carry_9_18), .ow_sum(w_sum_10_14), .ow_c(w_carry_10_14));
wire w_sum_10_12, w_carry_10_12;
math_adder_carry_save CSA_10_12(.i_a(w_carry_9_16), .i_b(w_carry_9_14), .i_c(w_carry_9_12), .ow_sum(w_sum_10_12), .ow_c(w_carry_10_12));
wire w_sum_10_10, w_carry_10_10;
math_adder_carry_save CSA_10_10(.i_a(w_carry_9_10), .i_b(w_carry_9_8), .i_c(w_carry_9_6), .ow_sum(w_sum_10_10), .ow_c(w_carry_10_10));
wire w_sum_10_8, w_carry_10_8;
math_adder_carry_save CSA_10_8(.i_a(w_carry_9_4), .i_b(w_carry_9_2), .i_c(w_sum_10_20), .ow_sum(w_sum_10_8), .ow_c(w_carry_10_8));
wire w_sum_10_6, w_carry_10_6;
math_adder_carry_save CSA_10_6(.i_a(w_sum_10_18), .i_b(w_sum_10_16), .i_c(w_sum_10_14), .ow_sum(w_sum_10_6), .ow_c(w_carry_10_6));
wire w_sum_10_4, w_carry_10_4;
math_adder_carry_save CSA_10_4(.i_a(w_sum_10_12), .i_b(w_sum_10_10), .i_c(w_sum_10_8), .ow_sum(w_sum_10_4), .ow_c(w_carry_10_4));
wire w_sum_10_2, w_carry_10_2;
math_adder_half HA_10_2(.i_a(w_sum_10_6), .i_b(w_sum_10_4), .ow_sum(w_sum_10_2), .ow_c(w_carry_10_2));
wire w_sum_11_22, w_carry_11_22;
math_adder_carry_save CSA_11_22(.i_a(w_pp_0_11), .i_b(w_pp_1_10), .i_c(w_pp_2_9), .ow_sum(w_sum_11_22), .ow_c(w_carry_11_22));
wire w_sum_11_20, w_carry_11_20;
math_adder_carry_save CSA_11_20(.i_a(w_pp_3_8), .i_b(w_pp_4_7), .i_c(w_pp_5_6), .ow_sum(w_sum_11_20), .ow_c(w_carry_11_20));
wire w_sum_11_18, w_carry_11_18;
math_adder_carry_save CSA_11_18(.i_a(w_pp_6_5), .i_b(w_pp_7_4), .i_c(w_pp_8_3), .ow_sum(w_sum_11_18), .ow_c(w_carry_11_18));
wire w_sum_11_16, w_carry_11_16;
math_adder_carry_save CSA_11_16(.i_a(w_pp_9_2), .i_b(w_pp_10_1), .i_c(w_pp_11_0), .ow_sum(w_sum_11_16), .ow_c(w_carry_11_16));
wire w_sum_11_14, w_carry_11_14;
math_adder_carry_save CSA_11_14(.i_a(w_carry_10_20), .i_b(w_carry_10_18), .i_c(w_carry_10_16), .ow_sum(w_sum_11_14), .ow_c(w_carry_11_14));
wire w_sum_11_12, w_carry_11_12;
math_adder_carry_save CSA_11_12(.i_a(w_carry_10_14), .i_b(w_carry_10_12), .i_c(w_carry_10_10), .ow_sum(w_sum_11_12), .ow_c(w_carry_11_12));
wire w_sum_11_10, w_carry_11_10;
math_adder_carry_save CSA_11_10(.i_a(w_carry_10_8), .i_b(w_carry_10_6), .i_c(w_carry_10_4), .ow_sum(w_sum_11_10), .ow_c(w_carry_11_10));
wire w_sum_11_8, w_carry_11_8;
math_adder_carry_save CSA_11_8(.i_a(w_carry_10_2), .i_b(w_sum_11_22), .i_c(w_sum_11_20), .ow_sum(w_sum_11_8), .ow_c(w_carry_11_8));
wire w_sum_11_6, w_carry_11_6;
math_adder_carry_save CSA_11_6(.i_a(w_sum_11_18), .i_b(w_sum_11_16), .i_c(w_sum_11_14), .ow_sum(w_sum_11_6), .ow_c(w_carry_11_6));
wire w_sum_11_4, w_carry_11_4;
math_adder_carry_save CSA_11_4(.i_a(w_sum_11_12), .i_b(w_sum_11_10), .i_c(w_sum_11_8), .ow_sum(w_sum_11_4), .ow_c(w_carry_11_4));
wire w_sum_11_2, w_carry_11_2;
math_adder_half HA_11_2(.i_a(w_sum_11_6), .i_b(w_sum_11_4), .ow_sum(w_sum_11_2), .ow_c(w_carry_11_2));
wire w_sum_12_24, w_carry_12_24;
math_adder_carry_save CSA_12_24(.i_a(w_pp_0_12), .i_b(w_pp_1_11), .i_c(w_pp_2_10), .ow_sum(w_sum_12_24), .ow_c(w_carry_12_24));
wire w_sum_12_22, w_carry_12_22;
math_adder_carry_save CSA_12_22(.i_a(w_pp_3_9), .i_b(w_pp_4_8), .i_c(w_pp_5_7), .ow_sum(w_sum_12_22), .ow_c(w_carry_12_22));
wire w_sum_12_20, w_carry_12_20;
math_adder_carry_save CSA_12_20(.i_a(w_pp_6_6), .i_b(w_pp_7_5), .i_c(w_pp_8_4), .ow_sum(w_sum_12_20), .ow_c(w_carry_12_20));
wire w_sum_12_18, w_carry_12_18;
math_adder_carry_save CSA_12_18(.i_a(w_pp_9_3), .i_b(w_pp_10_2), .i_c(w_pp_11_1), .ow_sum(w_sum_12_18), .ow_c(w_carry_12_18));
wire w_sum_12_16, w_carry_12_16;
math_adder_carry_save CSA_12_16(.i_a(w_pp_12_0), .i_b(w_carry_11_22), .i_c(w_carry_11_20), .ow_sum(w_sum_12_16), .ow_c(w_carry_12_16));
wire w_sum_12_14, w_carry_12_14;
math_adder_carry_save CSA_12_14(.i_a(w_carry_11_18), .i_b(w_carry_11_16), .i_c(w_carry_11_14), .ow_sum(w_sum_12_14), .ow_c(w_carry_12_14));
wire w_sum_12_12, w_carry_12_12;
math_adder_carry_save CSA_12_12(.i_a(w_carry_11_12), .i_b(w_carry_11_10), .i_c(w_carry_11_8), .ow_sum(w_sum_12_12), .ow_c(w_carry_12_12));
wire w_sum_12_10, w_carry_12_10;
math_adder_carry_save CSA_12_10(.i_a(w_carry_11_6), .i_b(w_carry_11_4), .i_c(w_carry_11_2), .ow_sum(w_sum_12_10), .ow_c(w_carry_12_10));
wire w_sum_12_8, w_carry_12_8;
math_adder_carry_save CSA_12_8(.i_a(w_sum_12_24), .i_b(w_sum_12_22), .i_c(w_sum_12_20), .ow_sum(w_sum_12_8), .ow_c(w_carry_12_8));
wire w_sum_12_6, w_carry_12_6;
math_adder_carry_save CSA_12_6(.i_a(w_sum_12_18), .i_b(w_sum_12_16), .i_c(w_sum_12_14), .ow_sum(w_sum_12_6), .ow_c(w_carry_12_6));
wire w_sum_12_4, w_carry_12_4;
math_adder_carry_save CSA_12_4(.i_a(w_sum_12_12), .i_b(w_sum_12_10), .i_c(w_sum_12_8), .ow_sum(w_sum_12_4), .ow_c(w_carry_12_4));
wire w_sum_12_2, w_carry_12_2;
math_adder_half HA_12_2(.i_a(w_sum_12_6), .i_b(w_sum_12_4), .ow_sum(w_sum_12_2), .ow_c(w_carry_12_2));
wire w_sum_13_26, w_carry_13_26;
math_adder_carry_save CSA_13_26(.i_a(w_pp_0_13), .i_b(w_pp_1_12), .i_c(w_pp_2_11), .ow_sum(w_sum_13_26), .ow_c(w_carry_13_26));
wire w_sum_13_24, w_carry_13_24;
math_adder_carry_save CSA_13_24(.i_a(w_pp_3_10), .i_b(w_pp_4_9), .i_c(w_pp_5_8), .ow_sum(w_sum_13_24), .ow_c(w_carry_13_24));
wire w_sum_13_22, w_carry_13_22;
math_adder_carry_save CSA_13_22(.i_a(w_pp_6_7), .i_b(w_pp_7_6), .i_c(w_pp_8_5), .ow_sum(w_sum_13_22), .ow_c(w_carry_13_22));
wire w_sum_13_20, w_carry_13_20;
math_adder_carry_save CSA_13_20(.i_a(w_pp_9_4), .i_b(w_pp_10_3), .i_c(w_pp_11_2), .ow_sum(w_sum_13_20), .ow_c(w_carry_13_20));
wire w_sum_13_18, w_carry_13_18;
math_adder_carry_save CSA_13_18(.i_a(w_pp_12_1), .i_b(w_pp_13_0), .i_c(w_carry_12_24), .ow_sum(w_sum_13_18), .ow_c(w_carry_13_18));
wire w_sum_13_16, w_carry_13_16;
math_adder_carry_save CSA_13_16(.i_a(w_carry_12_22), .i_b(w_carry_12_20), .i_c(w_carry_12_18), .ow_sum(w_sum_13_16), .ow_c(w_carry_13_16));
wire w_sum_13_14, w_carry_13_14;
math_adder_carry_save CSA_13_14(.i_a(w_carry_12_16), .i_b(w_carry_12_14), .i_c(w_carry_12_12), .ow_sum(w_sum_13_14), .ow_c(w_carry_13_14));
wire w_sum_13_12, w_carry_13_12;
math_adder_carry_save CSA_13_12(.i_a(w_carry_12_10), .i_b(w_carry_12_8), .i_c(w_carry_12_6), .ow_sum(w_sum_13_12), .ow_c(w_carry_13_12));
wire w_sum_13_10, w_carry_13_10;
math_adder_carry_save CSA_13_10(.i_a(w_carry_12_4), .i_b(w_carry_12_2), .i_c(w_sum_13_26), .ow_sum(w_sum_13_10), .ow_c(w_carry_13_10));
wire w_sum_13_8, w_carry_13_8;
math_adder_carry_save CSA_13_8(.i_a(w_sum_13_24), .i_b(w_sum_13_22), .i_c(w_sum_13_20), .ow_sum(w_sum_13_8), .ow_c(w_carry_13_8));
wire w_sum_13_6, w_carry_13_6;
math_adder_carry_save CSA_13_6(.i_a(w_sum_13_18), .i_b(w_sum_13_16), .i_c(w_sum_13_14), .ow_sum(w_sum_13_6), .ow_c(w_carry_13_6));
wire w_sum_13_4, w_carry_13_4;
math_adder_carry_save CSA_13_4(.i_a(w_sum_13_12), .i_b(w_sum_13_10), .i_c(w_sum_13_8), .ow_sum(w_sum_13_4), .ow_c(w_carry_13_4));
wire w_sum_13_2, w_carry_13_2;
math_adder_half HA_13_2(.i_a(w_sum_13_6), .i_b(w_sum_13_4), .ow_sum(w_sum_13_2), .ow_c(w_carry_13_2));
wire w_sum_14_28, w_carry_14_28;
math_adder_carry_save CSA_14_28(.i_a(w_pp_0_14), .i_b(w_pp_1_13), .i_c(w_pp_2_12), .ow_sum(w_sum_14_28), .ow_c(w_carry_14_28));
wire w_sum_14_26, w_carry_14_26;
math_adder_carry_save CSA_14_26(.i_a(w_pp_3_11), .i_b(w_pp_4_10), .i_c(w_pp_5_9), .ow_sum(w_sum_14_26), .ow_c(w_carry_14_26));
wire w_sum_14_24, w_carry_14_24;
math_adder_carry_save CSA_14_24(.i_a(w_pp_6_8), .i_b(w_pp_7_7), .i_c(w_pp_8_6), .ow_sum(w_sum_14_24), .ow_c(w_carry_14_24));
wire w_sum_14_22, w_carry_14_22;
math_adder_carry_save CSA_14_22(.i_a(w_pp_9_5), .i_b(w_pp_10_4), .i_c(w_pp_11_3), .ow_sum(w_sum_14_22), .ow_c(w_carry_14_22));
wire w_sum_14_20, w_carry_14_20;
math_adder_carry_save CSA_14_20(.i_a(w_pp_12_2), .i_b(w_pp_13_1), .i_c(w_pp_14_0), .ow_sum(w_sum_14_20), .ow_c(w_carry_14_20));
wire w_sum_14_18, w_carry_14_18;
math_adder_carry_save CSA_14_18(.i_a(w_carry_13_26), .i_b(w_carry_13_24), .i_c(w_carry_13_22), .ow_sum(w_sum_14_18), .ow_c(w_carry_14_18));
wire w_sum_14_16, w_carry_14_16;
math_adder_carry_save CSA_14_16(.i_a(w_carry_13_20), .i_b(w_carry_13_18), .i_c(w_carry_13_16), .ow_sum(w_sum_14_16), .ow_c(w_carry_14_16));
wire w_sum_14_14, w_carry_14_14;
math_adder_carry_save CSA_14_14(.i_a(w_carry_13_14), .i_b(w_carry_13_12), .i_c(w_carry_13_10), .ow_sum(w_sum_14_14), .ow_c(w_carry_14_14));
wire w_sum_14_12, w_carry_14_12;
math_adder_carry_save CSA_14_12(.i_a(w_carry_13_8), .i_b(w_carry_13_6), .i_c(w_carry_13_4), .ow_sum(w_sum_14_12), .ow_c(w_carry_14_12));
wire w_sum_14_10, w_carry_14_10;
math_adder_carry_save CSA_14_10(.i_a(w_carry_13_2), .i_b(w_sum_14_28), .i_c(w_sum_14_26), .ow_sum(w_sum_14_10), .ow_c(w_carry_14_10));
wire w_sum_14_8, w_carry_14_8;
math_adder_carry_save CSA_14_8(.i_a(w_sum_14_24), .i_b(w_sum_14_22), .i_c(w_sum_14_20), .ow_sum(w_sum_14_8), .ow_c(w_carry_14_8));
wire w_sum_14_6, w_carry_14_6;
math_adder_carry_save CSA_14_6(.i_a(w_sum_14_18), .i_b(w_sum_14_16), .i_c(w_sum_14_14), .ow_sum(w_sum_14_6), .ow_c(w_carry_14_6));
wire w_sum_14_4, w_carry_14_4;
math_adder_carry_save CSA_14_4(.i_a(w_sum_14_12), .i_b(w_sum_14_10), .i_c(w_sum_14_8), .ow_sum(w_sum_14_4), .ow_c(w_carry_14_4));
wire w_sum_14_2, w_carry_14_2;
math_adder_half HA_14_2(.i_a(w_sum_14_6), .i_b(w_sum_14_4), .ow_sum(w_sum_14_2), .ow_c(w_carry_14_2));
wire w_sum_15_30, w_carry_15_30;
math_adder_carry_save CSA_15_30(.i_a(w_pp_0_15), .i_b(w_pp_1_14), .i_c(w_pp_2_13), .ow_sum(w_sum_15_30), .ow_c(w_carry_15_30));
wire w_sum_15_28, w_carry_15_28;
math_adder_carry_save CSA_15_28(.i_a(w_pp_3_12), .i_b(w_pp_4_11), .i_c(w_pp_5_10), .ow_sum(w_sum_15_28), .ow_c(w_carry_15_28));
wire w_sum_15_26, w_carry_15_26;
math_adder_carry_save CSA_15_26(.i_a(w_pp_6_9), .i_b(w_pp_7_8), .i_c(w_pp_8_7), .ow_sum(w_sum_15_26), .ow_c(w_carry_15_26));
wire w_sum_15_24, w_carry_15_24;
math_adder_carry_save CSA_15_24(.i_a(w_pp_9_6), .i_b(w_pp_10_5), .i_c(w_pp_11_4), .ow_sum(w_sum_15_24), .ow_c(w_carry_15_24));
wire w_sum_15_22, w_carry_15_22;
math_adder_carry_save CSA_15_22(.i_a(w_pp_12_3), .i_b(w_pp_13_2), .i_c(w_pp_14_1), .ow_sum(w_sum_15_22), .ow_c(w_carry_15_22));
wire w_sum_15_20, w_carry_15_20;
math_adder_carry_save CSA_15_20(.i_a(w_pp_15_0), .i_b(w_carry_14_28), .i_c(w_carry_14_26), .ow_sum(w_sum_15_20), .ow_c(w_carry_15_20));
wire w_sum_15_18, w_carry_15_18;
math_adder_carry_save CSA_15_18(.i_a(w_carry_14_24), .i_b(w_carry_14_22), .i_c(w_carry_14_20), .ow_sum(w_sum_15_18), .ow_c(w_carry_15_18));
wire w_sum_15_16, w_carry_15_16;
math_adder_carry_save CSA_15_16(.i_a(w_carry_14_18), .i_b(w_carry_14_16), .i_c(w_carry_14_14), .ow_sum(w_sum_15_16), .ow_c(w_carry_15_16));
wire w_sum_15_14, w_carry_15_14;
math_adder_carry_save CSA_15_14(.i_a(w_carry_14_12), .i_b(w_carry_14_10), .i_c(w_carry_14_8), .ow_sum(w_sum_15_14), .ow_c(w_carry_15_14));
wire w_sum_15_12, w_carry_15_12;
math_adder_carry_save CSA_15_12(.i_a(w_carry_14_6), .i_b(w_carry_14_4), .i_c(w_carry_14_2), .ow_sum(w_sum_15_12), .ow_c(w_carry_15_12));
wire w_sum_15_10, w_carry_15_10;
math_adder_carry_save CSA_15_10(.i_a(w_sum_15_30), .i_b(w_sum_15_28), .i_c(w_sum_15_26), .ow_sum(w_sum_15_10), .ow_c(w_carry_15_10));
wire w_sum_15_8, w_carry_15_8;
math_adder_carry_save CSA_15_8(.i_a(w_sum_15_24), .i_b(w_sum_15_22), .i_c(w_sum_15_20), .ow_sum(w_sum_15_8), .ow_c(w_carry_15_8));
wire w_sum_15_6, w_carry_15_6;
math_adder_carry_save CSA_15_6(.i_a(w_sum_15_18), .i_b(w_sum_15_16), .i_c(w_sum_15_14), .ow_sum(w_sum_15_6), .ow_c(w_carry_15_6));
wire w_sum_15_4, w_carry_15_4;
math_adder_carry_save CSA_15_4(.i_a(w_sum_15_12), .i_b(w_sum_15_10), .i_c(w_sum_15_8), .ow_sum(w_sum_15_4), .ow_c(w_carry_15_4));
wire w_sum_15_2, w_carry_15_2;
math_adder_half HA_15_2(.i_a(w_sum_15_6), .i_b(w_sum_15_4), .ow_sum(w_sum_15_2), .ow_c(w_carry_15_2));
wire w_sum_16_32, w_carry_16_32;
math_adder_carry_save CSA_16_32(.i_a(w_pp_0_16), .i_b(w_pp_1_15), .i_c(w_pp_2_14), .ow_sum(w_sum_16_32), .ow_c(w_carry_16_32));
wire w_sum_16_30, w_carry_16_30;
math_adder_carry_save CSA_16_30(.i_a(w_pp_3_13), .i_b(w_pp_4_12), .i_c(w_pp_5_11), .ow_sum(w_sum_16_30), .ow_c(w_carry_16_30));
wire w_sum_16_28, w_carry_16_28;
math_adder_carry_save CSA_16_28(.i_a(w_pp_6_10), .i_b(w_pp_7_9), .i_c(w_pp_8_8), .ow_sum(w_sum_16_28), .ow_c(w_carry_16_28));
wire w_sum_16_26, w_carry_16_26;
math_adder_carry_save CSA_16_26(.i_a(w_pp_9_7), .i_b(w_pp_10_6), .i_c(w_pp_11_5), .ow_sum(w_sum_16_26), .ow_c(w_carry_16_26));
wire w_sum_16_24, w_carry_16_24;
math_adder_carry_save CSA_16_24(.i_a(w_pp_12_4), .i_b(w_pp_13_3), .i_c(w_pp_14_2), .ow_sum(w_sum_16_24), .ow_c(w_carry_16_24));
wire w_sum_16_22, w_carry_16_22;
math_adder_carry_save CSA_16_22(.i_a(w_pp_15_1), .i_b(w_pp_16_0), .i_c(w_carry_15_30), .ow_sum(w_sum_16_22), .ow_c(w_carry_16_22));
wire w_sum_16_20, w_carry_16_20;
math_adder_carry_save CSA_16_20(.i_a(w_carry_15_28), .i_b(w_carry_15_26), .i_c(w_carry_15_24), .ow_sum(w_sum_16_20), .ow_c(w_carry_16_20));
wire w_sum_16_18, w_carry_16_18;
math_adder_carry_save CSA_16_18(.i_a(w_carry_15_22), .i_b(w_carry_15_20), .i_c(w_carry_15_18), .ow_sum(w_sum_16_18), .ow_c(w_carry_16_18));
wire w_sum_16_16, w_carry_16_16;
math_adder_carry_save CSA_16_16(.i_a(w_carry_15_16), .i_b(w_carry_15_14), .i_c(w_carry_15_12), .ow_sum(w_sum_16_16), .ow_c(w_carry_16_16));
wire w_sum_16_14, w_carry_16_14;
math_adder_carry_save CSA_16_14(.i_a(w_carry_15_10), .i_b(w_carry_15_8), .i_c(w_carry_15_6), .ow_sum(w_sum_16_14), .ow_c(w_carry_16_14));
wire w_sum_16_12, w_carry_16_12;
math_adder_carry_save CSA_16_12(.i_a(w_carry_15_4), .i_b(w_carry_15_2), .i_c(w_sum_16_32), .ow_sum(w_sum_16_12), .ow_c(w_carry_16_12));
wire w_sum_16_10, w_carry_16_10;
math_adder_carry_save CSA_16_10(.i_a(w_sum_16_30), .i_b(w_sum_16_28), .i_c(w_sum_16_26), .ow_sum(w_sum_16_10), .ow_c(w_carry_16_10));
wire w_sum_16_8, w_carry_16_8;
math_adder_carry_save CSA_16_8(.i_a(w_sum_16_24), .i_b(w_sum_16_22), .i_c(w_sum_16_20), .ow_sum(w_sum_16_8), .ow_c(w_carry_16_8));
wire w_sum_16_6, w_carry_16_6;
math_adder_carry_save CSA_16_6(.i_a(w_sum_16_18), .i_b(w_sum_16_16), .i_c(w_sum_16_14), .ow_sum(w_sum_16_6), .ow_c(w_carry_16_6));
wire w_sum_16_4, w_carry_16_4;
math_adder_carry_save CSA_16_4(.i_a(w_sum_16_12), .i_b(w_sum_16_10), .i_c(w_sum_16_8), .ow_sum(w_sum_16_4), .ow_c(w_carry_16_4));
wire w_sum_16_2, w_carry_16_2;
math_adder_half HA_16_2(.i_a(w_sum_16_6), .i_b(w_sum_16_4), .ow_sum(w_sum_16_2), .ow_c(w_carry_16_2));
wire w_sum_17_34, w_carry_17_34;
math_adder_carry_save CSA_17_34(.i_a(w_pp_0_17), .i_b(w_pp_1_16), .i_c(w_pp_2_15), .ow_sum(w_sum_17_34), .ow_c(w_carry_17_34));
wire w_sum_17_32, w_carry_17_32;
math_adder_carry_save CSA_17_32(.i_a(w_pp_3_14), .i_b(w_pp_4_13), .i_c(w_pp_5_12), .ow_sum(w_sum_17_32), .ow_c(w_carry_17_32));
wire w_sum_17_30, w_carry_17_30;
math_adder_carry_save CSA_17_30(.i_a(w_pp_6_11), .i_b(w_pp_7_10), .i_c(w_pp_8_9), .ow_sum(w_sum_17_30), .ow_c(w_carry_17_30));
wire w_sum_17_28, w_carry_17_28;
math_adder_carry_save CSA_17_28(.i_a(w_pp_9_8), .i_b(w_pp_10_7), .i_c(w_pp_11_6), .ow_sum(w_sum_17_28), .ow_c(w_carry_17_28));
wire w_sum_17_26, w_carry_17_26;
math_adder_carry_save CSA_17_26(.i_a(w_pp_12_5), .i_b(w_pp_13_4), .i_c(w_pp_14_3), .ow_sum(w_sum_17_26), .ow_c(w_carry_17_26));
wire w_sum_17_24, w_carry_17_24;
math_adder_carry_save CSA_17_24(.i_a(w_pp_15_2), .i_b(w_pp_16_1), .i_c(w_pp_17_0), .ow_sum(w_sum_17_24), .ow_c(w_carry_17_24));
wire w_sum_17_22, w_carry_17_22;
math_adder_carry_save CSA_17_22(.i_a(w_carry_16_32), .i_b(w_carry_16_30), .i_c(w_carry_16_28), .ow_sum(w_sum_17_22), .ow_c(w_carry_17_22));
wire w_sum_17_20, w_carry_17_20;
math_adder_carry_save CSA_17_20(.i_a(w_carry_16_26), .i_b(w_carry_16_24), .i_c(w_carry_16_22), .ow_sum(w_sum_17_20), .ow_c(w_carry_17_20));
wire w_sum_17_18, w_carry_17_18;
math_adder_carry_save CSA_17_18(.i_a(w_carry_16_20), .i_b(w_carry_16_18), .i_c(w_carry_16_16), .ow_sum(w_sum_17_18), .ow_c(w_carry_17_18));
wire w_sum_17_16, w_carry_17_16;
math_adder_carry_save CSA_17_16(.i_a(w_carry_16_14), .i_b(w_carry_16_12), .i_c(w_carry_16_10), .ow_sum(w_sum_17_16), .ow_c(w_carry_17_16));
wire w_sum_17_14, w_carry_17_14;
math_adder_carry_save CSA_17_14(.i_a(w_carry_16_8), .i_b(w_carry_16_6), .i_c(w_carry_16_4), .ow_sum(w_sum_17_14), .ow_c(w_carry_17_14));
wire w_sum_17_12, w_carry_17_12;
math_adder_carry_save CSA_17_12(.i_a(w_carry_16_2), .i_b(w_sum_17_34), .i_c(w_sum_17_32), .ow_sum(w_sum_17_12), .ow_c(w_carry_17_12));
wire w_sum_17_10, w_carry_17_10;
math_adder_carry_save CSA_17_10(.i_a(w_sum_17_30), .i_b(w_sum_17_28), .i_c(w_sum_17_26), .ow_sum(w_sum_17_10), .ow_c(w_carry_17_10));
wire w_sum_17_8, w_carry_17_8;
math_adder_carry_save CSA_17_8(.i_a(w_sum_17_24), .i_b(w_sum_17_22), .i_c(w_sum_17_20), .ow_sum(w_sum_17_8), .ow_c(w_carry_17_8));
wire w_sum_17_6, w_carry_17_6;
math_adder_carry_save CSA_17_6(.i_a(w_sum_17_18), .i_b(w_sum_17_16), .i_c(w_sum_17_14), .ow_sum(w_sum_17_6), .ow_c(w_carry_17_6));
wire w_sum_17_4, w_carry_17_4;
math_adder_carry_save CSA_17_4(.i_a(w_sum_17_12), .i_b(w_sum_17_10), .i_c(w_sum_17_8), .ow_sum(w_sum_17_4), .ow_c(w_carry_17_4));
wire w_sum_17_2, w_carry_17_2;
math_adder_half HA_17_2(.i_a(w_sum_17_6), .i_b(w_sum_17_4), .ow_sum(w_sum_17_2), .ow_c(w_carry_17_2));
wire w_sum_18_36, w_carry_18_36;
math_adder_carry_save CSA_18_36(.i_a(w_pp_0_18), .i_b(w_pp_1_17), .i_c(w_pp_2_16), .ow_sum(w_sum_18_36), .ow_c(w_carry_18_36));
wire w_sum_18_34, w_carry_18_34;
math_adder_carry_save CSA_18_34(.i_a(w_pp_3_15), .i_b(w_pp_4_14), .i_c(w_pp_5_13), .ow_sum(w_sum_18_34), .ow_c(w_carry_18_34));
wire w_sum_18_32, w_carry_18_32;
math_adder_carry_save CSA_18_32(.i_a(w_pp_6_12), .i_b(w_pp_7_11), .i_c(w_pp_8_10), .ow_sum(w_sum_18_32), .ow_c(w_carry_18_32));
wire w_sum_18_30, w_carry_18_30;
math_adder_carry_save CSA_18_30(.i_a(w_pp_9_9), .i_b(w_pp_10_8), .i_c(w_pp_11_7), .ow_sum(w_sum_18_30), .ow_c(w_carry_18_30));
wire w_sum_18_28, w_carry_18_28;
math_adder_carry_save CSA_18_28(.i_a(w_pp_12_6), .i_b(w_pp_13_5), .i_c(w_pp_14_4), .ow_sum(w_sum_18_28), .ow_c(w_carry_18_28));
wire w_sum_18_26, w_carry_18_26;
math_adder_carry_save CSA_18_26(.i_a(w_pp_15_3), .i_b(w_pp_16_2), .i_c(w_pp_17_1), .ow_sum(w_sum_18_26), .ow_c(w_carry_18_26));
wire w_sum_18_24, w_carry_18_24;
math_adder_carry_save CSA_18_24(.i_a(w_pp_18_0), .i_b(w_carry_17_34), .i_c(w_carry_17_32), .ow_sum(w_sum_18_24), .ow_c(w_carry_18_24));
wire w_sum_18_22, w_carry_18_22;
math_adder_carry_save CSA_18_22(.i_a(w_carry_17_30), .i_b(w_carry_17_28), .i_c(w_carry_17_26), .ow_sum(w_sum_18_22), .ow_c(w_carry_18_22));
wire w_sum_18_20, w_carry_18_20;
math_adder_carry_save CSA_18_20(.i_a(w_carry_17_24), .i_b(w_carry_17_22), .i_c(w_carry_17_20), .ow_sum(w_sum_18_20), .ow_c(w_carry_18_20));
wire w_sum_18_18, w_carry_18_18;
math_adder_carry_save CSA_18_18(.i_a(w_carry_17_18), .i_b(w_carry_17_16), .i_c(w_carry_17_14), .ow_sum(w_sum_18_18), .ow_c(w_carry_18_18));
wire w_sum_18_16, w_carry_18_16;
math_adder_carry_save CSA_18_16(.i_a(w_carry_17_12), .i_b(w_carry_17_10), .i_c(w_carry_17_8), .ow_sum(w_sum_18_16), .ow_c(w_carry_18_16));
wire w_sum_18_14, w_carry_18_14;
math_adder_carry_save CSA_18_14(.i_a(w_carry_17_6), .i_b(w_carry_17_4), .i_c(w_carry_17_2), .ow_sum(w_sum_18_14), .ow_c(w_carry_18_14));
wire w_sum_18_12, w_carry_18_12;
math_adder_carry_save CSA_18_12(.i_a(w_sum_18_36), .i_b(w_sum_18_34), .i_c(w_sum_18_32), .ow_sum(w_sum_18_12), .ow_c(w_carry_18_12));
wire w_sum_18_10, w_carry_18_10;
math_adder_carry_save CSA_18_10(.i_a(w_sum_18_30), .i_b(w_sum_18_28), .i_c(w_sum_18_26), .ow_sum(w_sum_18_10), .ow_c(w_carry_18_10));
wire w_sum_18_8, w_carry_18_8;
math_adder_carry_save CSA_18_8(.i_a(w_sum_18_24), .i_b(w_sum_18_22), .i_c(w_sum_18_20), .ow_sum(w_sum_18_8), .ow_c(w_carry_18_8));
wire w_sum_18_6, w_carry_18_6;
math_adder_carry_save CSA_18_6(.i_a(w_sum_18_18), .i_b(w_sum_18_16), .i_c(w_sum_18_14), .ow_sum(w_sum_18_6), .ow_c(w_carry_18_6));
wire w_sum_18_4, w_carry_18_4;
math_adder_carry_save CSA_18_4(.i_a(w_sum_18_12), .i_b(w_sum_18_10), .i_c(w_sum_18_8), .ow_sum(w_sum_18_4), .ow_c(w_carry_18_4));
wire w_sum_18_2, w_carry_18_2;
math_adder_half HA_18_2(.i_a(w_sum_18_6), .i_b(w_sum_18_4), .ow_sum(w_sum_18_2), .ow_c(w_carry_18_2));
wire w_sum_19_38, w_carry_19_38;
math_adder_carry_save CSA_19_38(.i_a(w_pp_0_19), .i_b(w_pp_1_18), .i_c(w_pp_2_17), .ow_sum(w_sum_19_38), .ow_c(w_carry_19_38));
wire w_sum_19_36, w_carry_19_36;
math_adder_carry_save CSA_19_36(.i_a(w_pp_3_16), .i_b(w_pp_4_15), .i_c(w_pp_5_14), .ow_sum(w_sum_19_36), .ow_c(w_carry_19_36));
wire w_sum_19_34, w_carry_19_34;
math_adder_carry_save CSA_19_34(.i_a(w_pp_6_13), .i_b(w_pp_7_12), .i_c(w_pp_8_11), .ow_sum(w_sum_19_34), .ow_c(w_carry_19_34));
wire w_sum_19_32, w_carry_19_32;
math_adder_carry_save CSA_19_32(.i_a(w_pp_9_10), .i_b(w_pp_10_9), .i_c(w_pp_11_8), .ow_sum(w_sum_19_32), .ow_c(w_carry_19_32));
wire w_sum_19_30, w_carry_19_30;
math_adder_carry_save CSA_19_30(.i_a(w_pp_12_7), .i_b(w_pp_13_6), .i_c(w_pp_14_5), .ow_sum(w_sum_19_30), .ow_c(w_carry_19_30));
wire w_sum_19_28, w_carry_19_28;
math_adder_carry_save CSA_19_28(.i_a(w_pp_15_4), .i_b(w_pp_16_3), .i_c(w_pp_17_2), .ow_sum(w_sum_19_28), .ow_c(w_carry_19_28));
wire w_sum_19_26, w_carry_19_26;
math_adder_carry_save CSA_19_26(.i_a(w_pp_18_1), .i_b(w_pp_19_0), .i_c(w_carry_18_36), .ow_sum(w_sum_19_26), .ow_c(w_carry_19_26));
wire w_sum_19_24, w_carry_19_24;
math_adder_carry_save CSA_19_24(.i_a(w_carry_18_34), .i_b(w_carry_18_32), .i_c(w_carry_18_30), .ow_sum(w_sum_19_24), .ow_c(w_carry_19_24));
wire w_sum_19_22, w_carry_19_22;
math_adder_carry_save CSA_19_22(.i_a(w_carry_18_28), .i_b(w_carry_18_26), .i_c(w_carry_18_24), .ow_sum(w_sum_19_22), .ow_c(w_carry_19_22));
wire w_sum_19_20, w_carry_19_20;
math_adder_carry_save CSA_19_20(.i_a(w_carry_18_22), .i_b(w_carry_18_20), .i_c(w_carry_18_18), .ow_sum(w_sum_19_20), .ow_c(w_carry_19_20));
wire w_sum_19_18, w_carry_19_18;
math_adder_carry_save CSA_19_18(.i_a(w_carry_18_16), .i_b(w_carry_18_14), .i_c(w_carry_18_12), .ow_sum(w_sum_19_18), .ow_c(w_carry_19_18));
wire w_sum_19_16, w_carry_19_16;
math_adder_carry_save CSA_19_16(.i_a(w_carry_18_10), .i_b(w_carry_18_8), .i_c(w_carry_18_6), .ow_sum(w_sum_19_16), .ow_c(w_carry_19_16));
wire w_sum_19_14, w_carry_19_14;
math_adder_carry_save CSA_19_14(.i_a(w_carry_18_4), .i_b(w_carry_18_2), .i_c(w_sum_19_38), .ow_sum(w_sum_19_14), .ow_c(w_carry_19_14));
wire w_sum_19_12, w_carry_19_12;
math_adder_carry_save CSA_19_12(.i_a(w_sum_19_36), .i_b(w_sum_19_34), .i_c(w_sum_19_32), .ow_sum(w_sum_19_12), .ow_c(w_carry_19_12));
wire w_sum_19_10, w_carry_19_10;
math_adder_carry_save CSA_19_10(.i_a(w_sum_19_30), .i_b(w_sum_19_28), .i_c(w_sum_19_26), .ow_sum(w_sum_19_10), .ow_c(w_carry_19_10));
wire w_sum_19_8, w_carry_19_8;
math_adder_carry_save CSA_19_8(.i_a(w_sum_19_24), .i_b(w_sum_19_22), .i_c(w_sum_19_20), .ow_sum(w_sum_19_8), .ow_c(w_carry_19_8));
wire w_sum_19_6, w_carry_19_6;
math_adder_carry_save CSA_19_6(.i_a(w_sum_19_18), .i_b(w_sum_19_16), .i_c(w_sum_19_14), .ow_sum(w_sum_19_6), .ow_c(w_carry_19_6));
wire w_sum_19_4, w_carry_19_4;
math_adder_carry_save CSA_19_4(.i_a(w_sum_19_12), .i_b(w_sum_19_10), .i_c(w_sum_19_8), .ow_sum(w_sum_19_4), .ow_c(w_carry_19_4));
wire w_sum_19_2, w_carry_19_2;
math_adder_half HA_19_2(.i_a(w_sum_19_6), .i_b(w_sum_19_4), .ow_sum(w_sum_19_2), .ow_c(w_carry_19_2));
wire w_sum_20_40, w_carry_20_40;
math_adder_carry_save CSA_20_40(.i_a(w_pp_0_20), .i_b(w_pp_1_19), .i_c(w_pp_2_18), .ow_sum(w_sum_20_40), .ow_c(w_carry_20_40));
wire w_sum_20_38, w_carry_20_38;
math_adder_carry_save CSA_20_38(.i_a(w_pp_3_17), .i_b(w_pp_4_16), .i_c(w_pp_5_15), .ow_sum(w_sum_20_38), .ow_c(w_carry_20_38));
wire w_sum_20_36, w_carry_20_36;
math_adder_carry_save CSA_20_36(.i_a(w_pp_6_14), .i_b(w_pp_7_13), .i_c(w_pp_8_12), .ow_sum(w_sum_20_36), .ow_c(w_carry_20_36));
wire w_sum_20_34, w_carry_20_34;
math_adder_carry_save CSA_20_34(.i_a(w_pp_9_11), .i_b(w_pp_10_10), .i_c(w_pp_11_9), .ow_sum(w_sum_20_34), .ow_c(w_carry_20_34));
wire w_sum_20_32, w_carry_20_32;
math_adder_carry_save CSA_20_32(.i_a(w_pp_12_8), .i_b(w_pp_13_7), .i_c(w_pp_14_6), .ow_sum(w_sum_20_32), .ow_c(w_carry_20_32));
wire w_sum_20_30, w_carry_20_30;
math_adder_carry_save CSA_20_30(.i_a(w_pp_15_5), .i_b(w_pp_16_4), .i_c(w_pp_17_3), .ow_sum(w_sum_20_30), .ow_c(w_carry_20_30));
wire w_sum_20_28, w_carry_20_28;
math_adder_carry_save CSA_20_28(.i_a(w_pp_18_2), .i_b(w_pp_19_1), .i_c(w_pp_20_0), .ow_sum(w_sum_20_28), .ow_c(w_carry_20_28));
wire w_sum_20_26, w_carry_20_26;
math_adder_carry_save CSA_20_26(.i_a(w_carry_19_38), .i_b(w_carry_19_36), .i_c(w_carry_19_34), .ow_sum(w_sum_20_26), .ow_c(w_carry_20_26));
wire w_sum_20_24, w_carry_20_24;
math_adder_carry_save CSA_20_24(.i_a(w_carry_19_32), .i_b(w_carry_19_30), .i_c(w_carry_19_28), .ow_sum(w_sum_20_24), .ow_c(w_carry_20_24));
wire w_sum_20_22, w_carry_20_22;
math_adder_carry_save CSA_20_22(.i_a(w_carry_19_26), .i_b(w_carry_19_24), .i_c(w_carry_19_22), .ow_sum(w_sum_20_22), .ow_c(w_carry_20_22));
wire w_sum_20_20, w_carry_20_20;
math_adder_carry_save CSA_20_20(.i_a(w_carry_19_20), .i_b(w_carry_19_18), .i_c(w_carry_19_16), .ow_sum(w_sum_20_20), .ow_c(w_carry_20_20));
wire w_sum_20_18, w_carry_20_18;
math_adder_carry_save CSA_20_18(.i_a(w_carry_19_14), .i_b(w_carry_19_12), .i_c(w_carry_19_10), .ow_sum(w_sum_20_18), .ow_c(w_carry_20_18));
wire w_sum_20_16, w_carry_20_16;
math_adder_carry_save CSA_20_16(.i_a(w_carry_19_8), .i_b(w_carry_19_6), .i_c(w_carry_19_4), .ow_sum(w_sum_20_16), .ow_c(w_carry_20_16));
wire w_sum_20_14, w_carry_20_14;
math_adder_carry_save CSA_20_14(.i_a(w_carry_19_2), .i_b(w_sum_20_40), .i_c(w_sum_20_38), .ow_sum(w_sum_20_14), .ow_c(w_carry_20_14));
wire w_sum_20_12, w_carry_20_12;
math_adder_carry_save CSA_20_12(.i_a(w_sum_20_36), .i_b(w_sum_20_34), .i_c(w_sum_20_32), .ow_sum(w_sum_20_12), .ow_c(w_carry_20_12));
wire w_sum_20_10, w_carry_20_10;
math_adder_carry_save CSA_20_10(.i_a(w_sum_20_30), .i_b(w_sum_20_28), .i_c(w_sum_20_26), .ow_sum(w_sum_20_10), .ow_c(w_carry_20_10));
wire w_sum_20_8, w_carry_20_8;
math_adder_carry_save CSA_20_8(.i_a(w_sum_20_24), .i_b(w_sum_20_22), .i_c(w_sum_20_20), .ow_sum(w_sum_20_8), .ow_c(w_carry_20_8));
wire w_sum_20_6, w_carry_20_6;
math_adder_carry_save CSA_20_6(.i_a(w_sum_20_18), .i_b(w_sum_20_16), .i_c(w_sum_20_14), .ow_sum(w_sum_20_6), .ow_c(w_carry_20_6));
wire w_sum_20_4, w_carry_20_4;
math_adder_carry_save CSA_20_4(.i_a(w_sum_20_12), .i_b(w_sum_20_10), .i_c(w_sum_20_8), .ow_sum(w_sum_20_4), .ow_c(w_carry_20_4));
wire w_sum_20_2, w_carry_20_2;
math_adder_half HA_20_2(.i_a(w_sum_20_6), .i_b(w_sum_20_4), .ow_sum(w_sum_20_2), .ow_c(w_carry_20_2));
wire w_sum_21_42, w_carry_21_42;
math_adder_carry_save CSA_21_42(.i_a(w_pp_0_21), .i_b(w_pp_1_20), .i_c(w_pp_2_19), .ow_sum(w_sum_21_42), .ow_c(w_carry_21_42));
wire w_sum_21_40, w_carry_21_40;
math_adder_carry_save CSA_21_40(.i_a(w_pp_3_18), .i_b(w_pp_4_17), .i_c(w_pp_5_16), .ow_sum(w_sum_21_40), .ow_c(w_carry_21_40));
wire w_sum_21_38, w_carry_21_38;
math_adder_carry_save CSA_21_38(.i_a(w_pp_6_15), .i_b(w_pp_7_14), .i_c(w_pp_8_13), .ow_sum(w_sum_21_38), .ow_c(w_carry_21_38));
wire w_sum_21_36, w_carry_21_36;
math_adder_carry_save CSA_21_36(.i_a(w_pp_9_12), .i_b(w_pp_10_11), .i_c(w_pp_11_10), .ow_sum(w_sum_21_36), .ow_c(w_carry_21_36));
wire w_sum_21_34, w_carry_21_34;
math_adder_carry_save CSA_21_34(.i_a(w_pp_12_9), .i_b(w_pp_13_8), .i_c(w_pp_14_7), .ow_sum(w_sum_21_34), .ow_c(w_carry_21_34));
wire w_sum_21_32, w_carry_21_32;
math_adder_carry_save CSA_21_32(.i_a(w_pp_15_6), .i_b(w_pp_16_5), .i_c(w_pp_17_4), .ow_sum(w_sum_21_32), .ow_c(w_carry_21_32));
wire w_sum_21_30, w_carry_21_30;
math_adder_carry_save CSA_21_30(.i_a(w_pp_18_3), .i_b(w_pp_19_2), .i_c(w_pp_20_1), .ow_sum(w_sum_21_30), .ow_c(w_carry_21_30));
wire w_sum_21_28, w_carry_21_28;
math_adder_carry_save CSA_21_28(.i_a(w_pp_21_0), .i_b(w_carry_20_40), .i_c(w_carry_20_38), .ow_sum(w_sum_21_28), .ow_c(w_carry_21_28));
wire w_sum_21_26, w_carry_21_26;
math_adder_carry_save CSA_21_26(.i_a(w_carry_20_36), .i_b(w_carry_20_34), .i_c(w_carry_20_32), .ow_sum(w_sum_21_26), .ow_c(w_carry_21_26));
wire w_sum_21_24, w_carry_21_24;
math_adder_carry_save CSA_21_24(.i_a(w_carry_20_30), .i_b(w_carry_20_28), .i_c(w_carry_20_26), .ow_sum(w_sum_21_24), .ow_c(w_carry_21_24));
wire w_sum_21_22, w_carry_21_22;
math_adder_carry_save CSA_21_22(.i_a(w_carry_20_24), .i_b(w_carry_20_22), .i_c(w_carry_20_20), .ow_sum(w_sum_21_22), .ow_c(w_carry_21_22));
wire w_sum_21_20, w_carry_21_20;
math_adder_carry_save CSA_21_20(.i_a(w_carry_20_18), .i_b(w_carry_20_16), .i_c(w_carry_20_14), .ow_sum(w_sum_21_20), .ow_c(w_carry_21_20));
wire w_sum_21_18, w_carry_21_18;
math_adder_carry_save CSA_21_18(.i_a(w_carry_20_12), .i_b(w_carry_20_10), .i_c(w_carry_20_8), .ow_sum(w_sum_21_18), .ow_c(w_carry_21_18));
wire w_sum_21_16, w_carry_21_16;
math_adder_carry_save CSA_21_16(.i_a(w_carry_20_6), .i_b(w_carry_20_4), .i_c(w_carry_20_2), .ow_sum(w_sum_21_16), .ow_c(w_carry_21_16));
wire w_sum_21_14, w_carry_21_14;
math_adder_carry_save CSA_21_14(.i_a(w_sum_21_42), .i_b(w_sum_21_40), .i_c(w_sum_21_38), .ow_sum(w_sum_21_14), .ow_c(w_carry_21_14));
wire w_sum_21_12, w_carry_21_12;
math_adder_carry_save CSA_21_12(.i_a(w_sum_21_36), .i_b(w_sum_21_34), .i_c(w_sum_21_32), .ow_sum(w_sum_21_12), .ow_c(w_carry_21_12));
wire w_sum_21_10, w_carry_21_10;
math_adder_carry_save CSA_21_10(.i_a(w_sum_21_30), .i_b(w_sum_21_28), .i_c(w_sum_21_26), .ow_sum(w_sum_21_10), .ow_c(w_carry_21_10));
wire w_sum_21_8, w_carry_21_8;
math_adder_carry_save CSA_21_8(.i_a(w_sum_21_24), .i_b(w_sum_21_22), .i_c(w_sum_21_20), .ow_sum(w_sum_21_8), .ow_c(w_carry_21_8));
wire w_sum_21_6, w_carry_21_6;
math_adder_carry_save CSA_21_6(.i_a(w_sum_21_18), .i_b(w_sum_21_16), .i_c(w_sum_21_14), .ow_sum(w_sum_21_6), .ow_c(w_carry_21_6));
wire w_sum_21_4, w_carry_21_4;
math_adder_carry_save CSA_21_4(.i_a(w_sum_21_12), .i_b(w_sum_21_10), .i_c(w_sum_21_8), .ow_sum(w_sum_21_4), .ow_c(w_carry_21_4));
wire w_sum_21_2, w_carry_21_2;
math_adder_half HA_21_2(.i_a(w_sum_21_6), .i_b(w_sum_21_4), .ow_sum(w_sum_21_2), .ow_c(w_carry_21_2));
wire w_sum_22_44, w_carry_22_44;
math_adder_carry_save CSA_22_44(.i_a(w_pp_0_22), .i_b(w_pp_1_21), .i_c(w_pp_2_20), .ow_sum(w_sum_22_44), .ow_c(w_carry_22_44));
wire w_sum_22_42, w_carry_22_42;
math_adder_carry_save CSA_22_42(.i_a(w_pp_3_19), .i_b(w_pp_4_18), .i_c(w_pp_5_17), .ow_sum(w_sum_22_42), .ow_c(w_carry_22_42));
wire w_sum_22_40, w_carry_22_40;
math_adder_carry_save CSA_22_40(.i_a(w_pp_6_16), .i_b(w_pp_7_15), .i_c(w_pp_8_14), .ow_sum(w_sum_22_40), .ow_c(w_carry_22_40));
wire w_sum_22_38, w_carry_22_38;
math_adder_carry_save CSA_22_38(.i_a(w_pp_9_13), .i_b(w_pp_10_12), .i_c(w_pp_11_11), .ow_sum(w_sum_22_38), .ow_c(w_carry_22_38));
wire w_sum_22_36, w_carry_22_36;
math_adder_carry_save CSA_22_36(.i_a(w_pp_12_10), .i_b(w_pp_13_9), .i_c(w_pp_14_8), .ow_sum(w_sum_22_36), .ow_c(w_carry_22_36));
wire w_sum_22_34, w_carry_22_34;
math_adder_carry_save CSA_22_34(.i_a(w_pp_15_7), .i_b(w_pp_16_6), .i_c(w_pp_17_5), .ow_sum(w_sum_22_34), .ow_c(w_carry_22_34));
wire w_sum_22_32, w_carry_22_32;
math_adder_carry_save CSA_22_32(.i_a(w_pp_18_4), .i_b(w_pp_19_3), .i_c(w_pp_20_2), .ow_sum(w_sum_22_32), .ow_c(w_carry_22_32));
wire w_sum_22_30, w_carry_22_30;
math_adder_carry_save CSA_22_30(.i_a(w_pp_21_1), .i_b(w_pp_22_0), .i_c(w_carry_21_42), .ow_sum(w_sum_22_30), .ow_c(w_carry_22_30));
wire w_sum_22_28, w_carry_22_28;
math_adder_carry_save CSA_22_28(.i_a(w_carry_21_40), .i_b(w_carry_21_38), .i_c(w_carry_21_36), .ow_sum(w_sum_22_28), .ow_c(w_carry_22_28));
wire w_sum_22_26, w_carry_22_26;
math_adder_carry_save CSA_22_26(.i_a(w_carry_21_34), .i_b(w_carry_21_32), .i_c(w_carry_21_30), .ow_sum(w_sum_22_26), .ow_c(w_carry_22_26));
wire w_sum_22_24, w_carry_22_24;
math_adder_carry_save CSA_22_24(.i_a(w_carry_21_28), .i_b(w_carry_21_26), .i_c(w_carry_21_24), .ow_sum(w_sum_22_24), .ow_c(w_carry_22_24));
wire w_sum_22_22, w_carry_22_22;
math_adder_carry_save CSA_22_22(.i_a(w_carry_21_22), .i_b(w_carry_21_20), .i_c(w_carry_21_18), .ow_sum(w_sum_22_22), .ow_c(w_carry_22_22));
wire w_sum_22_20, w_carry_22_20;
math_adder_carry_save CSA_22_20(.i_a(w_carry_21_16), .i_b(w_carry_21_14), .i_c(w_carry_21_12), .ow_sum(w_sum_22_20), .ow_c(w_carry_22_20));
wire w_sum_22_18, w_carry_22_18;
math_adder_carry_save CSA_22_18(.i_a(w_carry_21_10), .i_b(w_carry_21_8), .i_c(w_carry_21_6), .ow_sum(w_sum_22_18), .ow_c(w_carry_22_18));
wire w_sum_22_16, w_carry_22_16;
math_adder_carry_save CSA_22_16(.i_a(w_carry_21_4), .i_b(w_carry_21_2), .i_c(w_sum_22_44), .ow_sum(w_sum_22_16), .ow_c(w_carry_22_16));
wire w_sum_22_14, w_carry_22_14;
math_adder_carry_save CSA_22_14(.i_a(w_sum_22_42), .i_b(w_sum_22_40), .i_c(w_sum_22_38), .ow_sum(w_sum_22_14), .ow_c(w_carry_22_14));
wire w_sum_22_12, w_carry_22_12;
math_adder_carry_save CSA_22_12(.i_a(w_sum_22_36), .i_b(w_sum_22_34), .i_c(w_sum_22_32), .ow_sum(w_sum_22_12), .ow_c(w_carry_22_12));
wire w_sum_22_10, w_carry_22_10;
math_adder_carry_save CSA_22_10(.i_a(w_sum_22_30), .i_b(w_sum_22_28), .i_c(w_sum_22_26), .ow_sum(w_sum_22_10), .ow_c(w_carry_22_10));
wire w_sum_22_8, w_carry_22_8;
math_adder_carry_save CSA_22_8(.i_a(w_sum_22_24), .i_b(w_sum_22_22), .i_c(w_sum_22_20), .ow_sum(w_sum_22_8), .ow_c(w_carry_22_8));
wire w_sum_22_6, w_carry_22_6;
math_adder_carry_save CSA_22_6(.i_a(w_sum_22_18), .i_b(w_sum_22_16), .i_c(w_sum_22_14), .ow_sum(w_sum_22_6), .ow_c(w_carry_22_6));
wire w_sum_22_4, w_carry_22_4;
math_adder_carry_save CSA_22_4(.i_a(w_sum_22_12), .i_b(w_sum_22_10), .i_c(w_sum_22_8), .ow_sum(w_sum_22_4), .ow_c(w_carry_22_4));
wire w_sum_22_2, w_carry_22_2;
math_adder_half HA_22_2(.i_a(w_sum_22_6), .i_b(w_sum_22_4), .ow_sum(w_sum_22_2), .ow_c(w_carry_22_2));
wire w_sum_23_46, w_carry_23_46;
math_adder_carry_save CSA_23_46(.i_a(w_pp_0_23), .i_b(w_pp_1_22), .i_c(w_pp_2_21), .ow_sum(w_sum_23_46), .ow_c(w_carry_23_46));
wire w_sum_23_44, w_carry_23_44;
math_adder_carry_save CSA_23_44(.i_a(w_pp_3_20), .i_b(w_pp_4_19), .i_c(w_pp_5_18), .ow_sum(w_sum_23_44), .ow_c(w_carry_23_44));
wire w_sum_23_42, w_carry_23_42;
math_adder_carry_save CSA_23_42(.i_a(w_pp_6_17), .i_b(w_pp_7_16), .i_c(w_pp_8_15), .ow_sum(w_sum_23_42), .ow_c(w_carry_23_42));
wire w_sum_23_40, w_carry_23_40;
math_adder_carry_save CSA_23_40(.i_a(w_pp_9_14), .i_b(w_pp_10_13), .i_c(w_pp_11_12), .ow_sum(w_sum_23_40), .ow_c(w_carry_23_40));
wire w_sum_23_38, w_carry_23_38;
math_adder_carry_save CSA_23_38(.i_a(w_pp_12_11), .i_b(w_pp_13_10), .i_c(w_pp_14_9), .ow_sum(w_sum_23_38), .ow_c(w_carry_23_38));
wire w_sum_23_36, w_carry_23_36;
math_adder_carry_save CSA_23_36(.i_a(w_pp_15_8), .i_b(w_pp_16_7), .i_c(w_pp_17_6), .ow_sum(w_sum_23_36), .ow_c(w_carry_23_36));
wire w_sum_23_34, w_carry_23_34;
math_adder_carry_save CSA_23_34(.i_a(w_pp_18_5), .i_b(w_pp_19_4), .i_c(w_pp_20_3), .ow_sum(w_sum_23_34), .ow_c(w_carry_23_34));
wire w_sum_23_32, w_carry_23_32;
math_adder_carry_save CSA_23_32(.i_a(w_pp_21_2), .i_b(w_pp_22_1), .i_c(w_pp_23_0), .ow_sum(w_sum_23_32), .ow_c(w_carry_23_32));
wire w_sum_23_30, w_carry_23_30;
math_adder_carry_save CSA_23_30(.i_a(w_carry_22_44), .i_b(w_carry_22_42), .i_c(w_carry_22_40), .ow_sum(w_sum_23_30), .ow_c(w_carry_23_30));
wire w_sum_23_28, w_carry_23_28;
math_adder_carry_save CSA_23_28(.i_a(w_carry_22_38), .i_b(w_carry_22_36), .i_c(w_carry_22_34), .ow_sum(w_sum_23_28), .ow_c(w_carry_23_28));
wire w_sum_23_26, w_carry_23_26;
math_adder_carry_save CSA_23_26(.i_a(w_carry_22_32), .i_b(w_carry_22_30), .i_c(w_carry_22_28), .ow_sum(w_sum_23_26), .ow_c(w_carry_23_26));
wire w_sum_23_24, w_carry_23_24;
math_adder_carry_save CSA_23_24(.i_a(w_carry_22_26), .i_b(w_carry_22_24), .i_c(w_carry_22_22), .ow_sum(w_sum_23_24), .ow_c(w_carry_23_24));
wire w_sum_23_22, w_carry_23_22;
math_adder_carry_save CSA_23_22(.i_a(w_carry_22_20), .i_b(w_carry_22_18), .i_c(w_carry_22_16), .ow_sum(w_sum_23_22), .ow_c(w_carry_23_22));
wire w_sum_23_20, w_carry_23_20;
math_adder_carry_save CSA_23_20(.i_a(w_carry_22_14), .i_b(w_carry_22_12), .i_c(w_carry_22_10), .ow_sum(w_sum_23_20), .ow_c(w_carry_23_20));
wire w_sum_23_18, w_carry_23_18;
math_adder_carry_save CSA_23_18(.i_a(w_carry_22_8), .i_b(w_carry_22_6), .i_c(w_carry_22_4), .ow_sum(w_sum_23_18), .ow_c(w_carry_23_18));
wire w_sum_23_16, w_carry_23_16;
math_adder_carry_save CSA_23_16(.i_a(w_carry_22_2), .i_b(w_sum_23_46), .i_c(w_sum_23_44), .ow_sum(w_sum_23_16), .ow_c(w_carry_23_16));
wire w_sum_23_14, w_carry_23_14;
math_adder_carry_save CSA_23_14(.i_a(w_sum_23_42), .i_b(w_sum_23_40), .i_c(w_sum_23_38), .ow_sum(w_sum_23_14), .ow_c(w_carry_23_14));
wire w_sum_23_12, w_carry_23_12;
math_adder_carry_save CSA_23_12(.i_a(w_sum_23_36), .i_b(w_sum_23_34), .i_c(w_sum_23_32), .ow_sum(w_sum_23_12), .ow_c(w_carry_23_12));
wire w_sum_23_10, w_carry_23_10;
math_adder_carry_save CSA_23_10(.i_a(w_sum_23_30), .i_b(w_sum_23_28), .i_c(w_sum_23_26), .ow_sum(w_sum_23_10), .ow_c(w_carry_23_10));
wire w_sum_23_8, w_carry_23_8;
math_adder_carry_save CSA_23_8(.i_a(w_sum_23_24), .i_b(w_sum_23_22), .i_c(w_sum_23_20), .ow_sum(w_sum_23_8), .ow_c(w_carry_23_8));
wire w_sum_23_6, w_carry_23_6;
math_adder_carry_save CSA_23_6(.i_a(w_sum_23_18), .i_b(w_sum_23_16), .i_c(w_sum_23_14), .ow_sum(w_sum_23_6), .ow_c(w_carry_23_6));
wire w_sum_23_4, w_carry_23_4;
math_adder_carry_save CSA_23_4(.i_a(w_sum_23_12), .i_b(w_sum_23_10), .i_c(w_sum_23_8), .ow_sum(w_sum_23_4), .ow_c(w_carry_23_4));
wire w_sum_23_2, w_carry_23_2;
math_adder_half HA_23_2(.i_a(w_sum_23_6), .i_b(w_sum_23_4), .ow_sum(w_sum_23_2), .ow_c(w_carry_23_2));
wire w_sum_24_48, w_carry_24_48;
math_adder_carry_save CSA_24_48(.i_a(w_pp_0_24), .i_b(w_pp_1_23), .i_c(w_pp_2_22), .ow_sum(w_sum_24_48), .ow_c(w_carry_24_48));
wire w_sum_24_46, w_carry_24_46;
math_adder_carry_save CSA_24_46(.i_a(w_pp_3_21), .i_b(w_pp_4_20), .i_c(w_pp_5_19), .ow_sum(w_sum_24_46), .ow_c(w_carry_24_46));
wire w_sum_24_44, w_carry_24_44;
math_adder_carry_save CSA_24_44(.i_a(w_pp_6_18), .i_b(w_pp_7_17), .i_c(w_pp_8_16), .ow_sum(w_sum_24_44), .ow_c(w_carry_24_44));
wire w_sum_24_42, w_carry_24_42;
math_adder_carry_save CSA_24_42(.i_a(w_pp_9_15), .i_b(w_pp_10_14), .i_c(w_pp_11_13), .ow_sum(w_sum_24_42), .ow_c(w_carry_24_42));
wire w_sum_24_40, w_carry_24_40;
math_adder_carry_save CSA_24_40(.i_a(w_pp_12_12), .i_b(w_pp_13_11), .i_c(w_pp_14_10), .ow_sum(w_sum_24_40), .ow_c(w_carry_24_40));
wire w_sum_24_38, w_carry_24_38;
math_adder_carry_save CSA_24_38(.i_a(w_pp_15_9), .i_b(w_pp_16_8), .i_c(w_pp_17_7), .ow_sum(w_sum_24_38), .ow_c(w_carry_24_38));
wire w_sum_24_36, w_carry_24_36;
math_adder_carry_save CSA_24_36(.i_a(w_pp_18_6), .i_b(w_pp_19_5), .i_c(w_pp_20_4), .ow_sum(w_sum_24_36), .ow_c(w_carry_24_36));
wire w_sum_24_34, w_carry_24_34;
math_adder_carry_save CSA_24_34(.i_a(w_pp_21_3), .i_b(w_pp_22_2), .i_c(w_pp_23_1), .ow_sum(w_sum_24_34), .ow_c(w_carry_24_34));
wire w_sum_24_32, w_carry_24_32;
math_adder_carry_save CSA_24_32(.i_a(w_pp_24_0), .i_b(w_carry_23_46), .i_c(w_carry_23_44), .ow_sum(w_sum_24_32), .ow_c(w_carry_24_32));
wire w_sum_24_30, w_carry_24_30;
math_adder_carry_save CSA_24_30(.i_a(w_carry_23_42), .i_b(w_carry_23_40), .i_c(w_carry_23_38), .ow_sum(w_sum_24_30), .ow_c(w_carry_24_30));
wire w_sum_24_28, w_carry_24_28;
math_adder_carry_save CSA_24_28(.i_a(w_carry_23_36), .i_b(w_carry_23_34), .i_c(w_carry_23_32), .ow_sum(w_sum_24_28), .ow_c(w_carry_24_28));
wire w_sum_24_26, w_carry_24_26;
math_adder_carry_save CSA_24_26(.i_a(w_carry_23_30), .i_b(w_carry_23_28), .i_c(w_carry_23_26), .ow_sum(w_sum_24_26), .ow_c(w_carry_24_26));
wire w_sum_24_24, w_carry_24_24;
math_adder_carry_save CSA_24_24(.i_a(w_carry_23_24), .i_b(w_carry_23_22), .i_c(w_carry_23_20), .ow_sum(w_sum_24_24), .ow_c(w_carry_24_24));
wire w_sum_24_22, w_carry_24_22;
math_adder_carry_save CSA_24_22(.i_a(w_carry_23_18), .i_b(w_carry_23_16), .i_c(w_carry_23_14), .ow_sum(w_sum_24_22), .ow_c(w_carry_24_22));
wire w_sum_24_20, w_carry_24_20;
math_adder_carry_save CSA_24_20(.i_a(w_carry_23_12), .i_b(w_carry_23_10), .i_c(w_carry_23_8), .ow_sum(w_sum_24_20), .ow_c(w_carry_24_20));
wire w_sum_24_18, w_carry_24_18;
math_adder_carry_save CSA_24_18(.i_a(w_carry_23_6), .i_b(w_carry_23_4), .i_c(w_carry_23_2), .ow_sum(w_sum_24_18), .ow_c(w_carry_24_18));
wire w_sum_24_16, w_carry_24_16;
math_adder_carry_save CSA_24_16(.i_a(w_sum_24_48), .i_b(w_sum_24_46), .i_c(w_sum_24_44), .ow_sum(w_sum_24_16), .ow_c(w_carry_24_16));
wire w_sum_24_14, w_carry_24_14;
math_adder_carry_save CSA_24_14(.i_a(w_sum_24_42), .i_b(w_sum_24_40), .i_c(w_sum_24_38), .ow_sum(w_sum_24_14), .ow_c(w_carry_24_14));
wire w_sum_24_12, w_carry_24_12;
math_adder_carry_save CSA_24_12(.i_a(w_sum_24_36), .i_b(w_sum_24_34), .i_c(w_sum_24_32), .ow_sum(w_sum_24_12), .ow_c(w_carry_24_12));
wire w_sum_24_10, w_carry_24_10;
math_adder_carry_save CSA_24_10(.i_a(w_sum_24_30), .i_b(w_sum_24_28), .i_c(w_sum_24_26), .ow_sum(w_sum_24_10), .ow_c(w_carry_24_10));
wire w_sum_24_8, w_carry_24_8;
math_adder_carry_save CSA_24_8(.i_a(w_sum_24_24), .i_b(w_sum_24_22), .i_c(w_sum_24_20), .ow_sum(w_sum_24_8), .ow_c(w_carry_24_8));
wire w_sum_24_6, w_carry_24_6;
math_adder_carry_save CSA_24_6(.i_a(w_sum_24_18), .i_b(w_sum_24_16), .i_c(w_sum_24_14), .ow_sum(w_sum_24_6), .ow_c(w_carry_24_6));
wire w_sum_24_4, w_carry_24_4;
math_adder_carry_save CSA_24_4(.i_a(w_sum_24_12), .i_b(w_sum_24_10), .i_c(w_sum_24_8), .ow_sum(w_sum_24_4), .ow_c(w_carry_24_4));
wire w_sum_24_2, w_carry_24_2;
math_adder_half HA_24_2(.i_a(w_sum_24_6), .i_b(w_sum_24_4), .ow_sum(w_sum_24_2), .ow_c(w_carry_24_2));
wire w_sum_25_50, w_carry_25_50;
math_adder_carry_save CSA_25_50(.i_a(w_pp_0_25), .i_b(w_pp_1_24), .i_c(w_pp_2_23), .ow_sum(w_sum_25_50), .ow_c(w_carry_25_50));
wire w_sum_25_48, w_carry_25_48;
math_adder_carry_save CSA_25_48(.i_a(w_pp_3_22), .i_b(w_pp_4_21), .i_c(w_pp_5_20), .ow_sum(w_sum_25_48), .ow_c(w_carry_25_48));
wire w_sum_25_46, w_carry_25_46;
math_adder_carry_save CSA_25_46(.i_a(w_pp_6_19), .i_b(w_pp_7_18), .i_c(w_pp_8_17), .ow_sum(w_sum_25_46), .ow_c(w_carry_25_46));
wire w_sum_25_44, w_carry_25_44;
math_adder_carry_save CSA_25_44(.i_a(w_pp_9_16), .i_b(w_pp_10_15), .i_c(w_pp_11_14), .ow_sum(w_sum_25_44), .ow_c(w_carry_25_44));
wire w_sum_25_42, w_carry_25_42;
math_adder_carry_save CSA_25_42(.i_a(w_pp_12_13), .i_b(w_pp_13_12), .i_c(w_pp_14_11), .ow_sum(w_sum_25_42), .ow_c(w_carry_25_42));
wire w_sum_25_40, w_carry_25_40;
math_adder_carry_save CSA_25_40(.i_a(w_pp_15_10), .i_b(w_pp_16_9), .i_c(w_pp_17_8), .ow_sum(w_sum_25_40), .ow_c(w_carry_25_40));
wire w_sum_25_38, w_carry_25_38;
math_adder_carry_save CSA_25_38(.i_a(w_pp_18_7), .i_b(w_pp_19_6), .i_c(w_pp_20_5), .ow_sum(w_sum_25_38), .ow_c(w_carry_25_38));
wire w_sum_25_36, w_carry_25_36;
math_adder_carry_save CSA_25_36(.i_a(w_pp_21_4), .i_b(w_pp_22_3), .i_c(w_pp_23_2), .ow_sum(w_sum_25_36), .ow_c(w_carry_25_36));
wire w_sum_25_34, w_carry_25_34;
math_adder_carry_save CSA_25_34(.i_a(w_pp_24_1), .i_b(w_pp_25_0), .i_c(w_carry_24_48), .ow_sum(w_sum_25_34), .ow_c(w_carry_25_34));
wire w_sum_25_32, w_carry_25_32;
math_adder_carry_save CSA_25_32(.i_a(w_carry_24_46), .i_b(w_carry_24_44), .i_c(w_carry_24_42), .ow_sum(w_sum_25_32), .ow_c(w_carry_25_32));
wire w_sum_25_30, w_carry_25_30;
math_adder_carry_save CSA_25_30(.i_a(w_carry_24_40), .i_b(w_carry_24_38), .i_c(w_carry_24_36), .ow_sum(w_sum_25_30), .ow_c(w_carry_25_30));
wire w_sum_25_28, w_carry_25_28;
math_adder_carry_save CSA_25_28(.i_a(w_carry_24_34), .i_b(w_carry_24_32), .i_c(w_carry_24_30), .ow_sum(w_sum_25_28), .ow_c(w_carry_25_28));
wire w_sum_25_26, w_carry_25_26;
math_adder_carry_save CSA_25_26(.i_a(w_carry_24_28), .i_b(w_carry_24_26), .i_c(w_carry_24_24), .ow_sum(w_sum_25_26), .ow_c(w_carry_25_26));
wire w_sum_25_24, w_carry_25_24;
math_adder_carry_save CSA_25_24(.i_a(w_carry_24_22), .i_b(w_carry_24_20), .i_c(w_carry_24_18), .ow_sum(w_sum_25_24), .ow_c(w_carry_25_24));
wire w_sum_25_22, w_carry_25_22;
math_adder_carry_save CSA_25_22(.i_a(w_carry_24_16), .i_b(w_carry_24_14), .i_c(w_carry_24_12), .ow_sum(w_sum_25_22), .ow_c(w_carry_25_22));
wire w_sum_25_20, w_carry_25_20;
math_adder_carry_save CSA_25_20(.i_a(w_carry_24_10), .i_b(w_carry_24_8), .i_c(w_carry_24_6), .ow_sum(w_sum_25_20), .ow_c(w_carry_25_20));
wire w_sum_25_18, w_carry_25_18;
math_adder_carry_save CSA_25_18(.i_a(w_carry_24_4), .i_b(w_carry_24_2), .i_c(w_sum_25_50), .ow_sum(w_sum_25_18), .ow_c(w_carry_25_18));
wire w_sum_25_16, w_carry_25_16;
math_adder_carry_save CSA_25_16(.i_a(w_sum_25_48), .i_b(w_sum_25_46), .i_c(w_sum_25_44), .ow_sum(w_sum_25_16), .ow_c(w_carry_25_16));
wire w_sum_25_14, w_carry_25_14;
math_adder_carry_save CSA_25_14(.i_a(w_sum_25_42), .i_b(w_sum_25_40), .i_c(w_sum_25_38), .ow_sum(w_sum_25_14), .ow_c(w_carry_25_14));
wire w_sum_25_12, w_carry_25_12;
math_adder_carry_save CSA_25_12(.i_a(w_sum_25_36), .i_b(w_sum_25_34), .i_c(w_sum_25_32), .ow_sum(w_sum_25_12), .ow_c(w_carry_25_12));
wire w_sum_25_10, w_carry_25_10;
math_adder_carry_save CSA_25_10(.i_a(w_sum_25_30), .i_b(w_sum_25_28), .i_c(w_sum_25_26), .ow_sum(w_sum_25_10), .ow_c(w_carry_25_10));
wire w_sum_25_8, w_carry_25_8;
math_adder_carry_save CSA_25_8(.i_a(w_sum_25_24), .i_b(w_sum_25_22), .i_c(w_sum_25_20), .ow_sum(w_sum_25_8), .ow_c(w_carry_25_8));
wire w_sum_25_6, w_carry_25_6;
math_adder_carry_save CSA_25_6(.i_a(w_sum_25_18), .i_b(w_sum_25_16), .i_c(w_sum_25_14), .ow_sum(w_sum_25_6), .ow_c(w_carry_25_6));
wire w_sum_25_4, w_carry_25_4;
math_adder_carry_save CSA_25_4(.i_a(w_sum_25_12), .i_b(w_sum_25_10), .i_c(w_sum_25_8), .ow_sum(w_sum_25_4), .ow_c(w_carry_25_4));
wire w_sum_25_2, w_carry_25_2;
math_adder_half HA_25_2(.i_a(w_sum_25_6), .i_b(w_sum_25_4), .ow_sum(w_sum_25_2), .ow_c(w_carry_25_2));
wire w_sum_26_52, w_carry_26_52;
math_adder_carry_save CSA_26_52(.i_a(w_pp_0_26), .i_b(w_pp_1_25), .i_c(w_pp_2_24), .ow_sum(w_sum_26_52), .ow_c(w_carry_26_52));
wire w_sum_26_50, w_carry_26_50;
math_adder_carry_save CSA_26_50(.i_a(w_pp_3_23), .i_b(w_pp_4_22), .i_c(w_pp_5_21), .ow_sum(w_sum_26_50), .ow_c(w_carry_26_50));
wire w_sum_26_48, w_carry_26_48;
math_adder_carry_save CSA_26_48(.i_a(w_pp_6_20), .i_b(w_pp_7_19), .i_c(w_pp_8_18), .ow_sum(w_sum_26_48), .ow_c(w_carry_26_48));
wire w_sum_26_46, w_carry_26_46;
math_adder_carry_save CSA_26_46(.i_a(w_pp_9_17), .i_b(w_pp_10_16), .i_c(w_pp_11_15), .ow_sum(w_sum_26_46), .ow_c(w_carry_26_46));
wire w_sum_26_44, w_carry_26_44;
math_adder_carry_save CSA_26_44(.i_a(w_pp_12_14), .i_b(w_pp_13_13), .i_c(w_pp_14_12), .ow_sum(w_sum_26_44), .ow_c(w_carry_26_44));
wire w_sum_26_42, w_carry_26_42;
math_adder_carry_save CSA_26_42(.i_a(w_pp_15_11), .i_b(w_pp_16_10), .i_c(w_pp_17_9), .ow_sum(w_sum_26_42), .ow_c(w_carry_26_42));
wire w_sum_26_40, w_carry_26_40;
math_adder_carry_save CSA_26_40(.i_a(w_pp_18_8), .i_b(w_pp_19_7), .i_c(w_pp_20_6), .ow_sum(w_sum_26_40), .ow_c(w_carry_26_40));
wire w_sum_26_38, w_carry_26_38;
math_adder_carry_save CSA_26_38(.i_a(w_pp_21_5), .i_b(w_pp_22_4), .i_c(w_pp_23_3), .ow_sum(w_sum_26_38), .ow_c(w_carry_26_38));
wire w_sum_26_36, w_carry_26_36;
math_adder_carry_save CSA_26_36(.i_a(w_pp_24_2), .i_b(w_pp_25_1), .i_c(w_pp_26_0), .ow_sum(w_sum_26_36), .ow_c(w_carry_26_36));
wire w_sum_26_34, w_carry_26_34;
math_adder_carry_save CSA_26_34(.i_a(w_carry_25_50), .i_b(w_carry_25_48), .i_c(w_carry_25_46), .ow_sum(w_sum_26_34), .ow_c(w_carry_26_34));
wire w_sum_26_32, w_carry_26_32;
math_adder_carry_save CSA_26_32(.i_a(w_carry_25_44), .i_b(w_carry_25_42), .i_c(w_carry_25_40), .ow_sum(w_sum_26_32), .ow_c(w_carry_26_32));
wire w_sum_26_30, w_carry_26_30;
math_adder_carry_save CSA_26_30(.i_a(w_carry_25_38), .i_b(w_carry_25_36), .i_c(w_carry_25_34), .ow_sum(w_sum_26_30), .ow_c(w_carry_26_30));
wire w_sum_26_28, w_carry_26_28;
math_adder_carry_save CSA_26_28(.i_a(w_carry_25_32), .i_b(w_carry_25_30), .i_c(w_carry_25_28), .ow_sum(w_sum_26_28), .ow_c(w_carry_26_28));
wire w_sum_26_26, w_carry_26_26;
math_adder_carry_save CSA_26_26(.i_a(w_carry_25_26), .i_b(w_carry_25_24), .i_c(w_carry_25_22), .ow_sum(w_sum_26_26), .ow_c(w_carry_26_26));
wire w_sum_26_24, w_carry_26_24;
math_adder_carry_save CSA_26_24(.i_a(w_carry_25_20), .i_b(w_carry_25_18), .i_c(w_carry_25_16), .ow_sum(w_sum_26_24), .ow_c(w_carry_26_24));
wire w_sum_26_22, w_carry_26_22;
math_adder_carry_save CSA_26_22(.i_a(w_carry_25_14), .i_b(w_carry_25_12), .i_c(w_carry_25_10), .ow_sum(w_sum_26_22), .ow_c(w_carry_26_22));
wire w_sum_26_20, w_carry_26_20;
math_adder_carry_save CSA_26_20(.i_a(w_carry_25_8), .i_b(w_carry_25_6), .i_c(w_carry_25_4), .ow_sum(w_sum_26_20), .ow_c(w_carry_26_20));
wire w_sum_26_18, w_carry_26_18;
math_adder_carry_save CSA_26_18(.i_a(w_carry_25_2), .i_b(w_sum_26_52), .i_c(w_sum_26_50), .ow_sum(w_sum_26_18), .ow_c(w_carry_26_18));
wire w_sum_26_16, w_carry_26_16;
math_adder_carry_save CSA_26_16(.i_a(w_sum_26_48), .i_b(w_sum_26_46), .i_c(w_sum_26_44), .ow_sum(w_sum_26_16), .ow_c(w_carry_26_16));
wire w_sum_26_14, w_carry_26_14;
math_adder_carry_save CSA_26_14(.i_a(w_sum_26_42), .i_b(w_sum_26_40), .i_c(w_sum_26_38), .ow_sum(w_sum_26_14), .ow_c(w_carry_26_14));
wire w_sum_26_12, w_carry_26_12;
math_adder_carry_save CSA_26_12(.i_a(w_sum_26_36), .i_b(w_sum_26_34), .i_c(w_sum_26_32), .ow_sum(w_sum_26_12), .ow_c(w_carry_26_12));
wire w_sum_26_10, w_carry_26_10;
math_adder_carry_save CSA_26_10(.i_a(w_sum_26_30), .i_b(w_sum_26_28), .i_c(w_sum_26_26), .ow_sum(w_sum_26_10), .ow_c(w_carry_26_10));
wire w_sum_26_8, w_carry_26_8;
math_adder_carry_save CSA_26_8(.i_a(w_sum_26_24), .i_b(w_sum_26_22), .i_c(w_sum_26_20), .ow_sum(w_sum_26_8), .ow_c(w_carry_26_8));
wire w_sum_26_6, w_carry_26_6;
math_adder_carry_save CSA_26_6(.i_a(w_sum_26_18), .i_b(w_sum_26_16), .i_c(w_sum_26_14), .ow_sum(w_sum_26_6), .ow_c(w_carry_26_6));
wire w_sum_26_4, w_carry_26_4;
math_adder_carry_save CSA_26_4(.i_a(w_sum_26_12), .i_b(w_sum_26_10), .i_c(w_sum_26_8), .ow_sum(w_sum_26_4), .ow_c(w_carry_26_4));
wire w_sum_26_2, w_carry_26_2;
math_adder_half HA_26_2(.i_a(w_sum_26_6), .i_b(w_sum_26_4), .ow_sum(w_sum_26_2), .ow_c(w_carry_26_2));
wire w_sum_27_54, w_carry_27_54;
math_adder_carry_save CSA_27_54(.i_a(w_pp_0_27), .i_b(w_pp_1_26), .i_c(w_pp_2_25), .ow_sum(w_sum_27_54), .ow_c(w_carry_27_54));
wire w_sum_27_52, w_carry_27_52;
math_adder_carry_save CSA_27_52(.i_a(w_pp_3_24), .i_b(w_pp_4_23), .i_c(w_pp_5_22), .ow_sum(w_sum_27_52), .ow_c(w_carry_27_52));
wire w_sum_27_50, w_carry_27_50;
math_adder_carry_save CSA_27_50(.i_a(w_pp_6_21), .i_b(w_pp_7_20), .i_c(w_pp_8_19), .ow_sum(w_sum_27_50), .ow_c(w_carry_27_50));
wire w_sum_27_48, w_carry_27_48;
math_adder_carry_save CSA_27_48(.i_a(w_pp_9_18), .i_b(w_pp_10_17), .i_c(w_pp_11_16), .ow_sum(w_sum_27_48), .ow_c(w_carry_27_48));
wire w_sum_27_46, w_carry_27_46;
math_adder_carry_save CSA_27_46(.i_a(w_pp_12_15), .i_b(w_pp_13_14), .i_c(w_pp_14_13), .ow_sum(w_sum_27_46), .ow_c(w_carry_27_46));
wire w_sum_27_44, w_carry_27_44;
math_adder_carry_save CSA_27_44(.i_a(w_pp_15_12), .i_b(w_pp_16_11), .i_c(w_pp_17_10), .ow_sum(w_sum_27_44), .ow_c(w_carry_27_44));
wire w_sum_27_42, w_carry_27_42;
math_adder_carry_save CSA_27_42(.i_a(w_pp_18_9), .i_b(w_pp_19_8), .i_c(w_pp_20_7), .ow_sum(w_sum_27_42), .ow_c(w_carry_27_42));
wire w_sum_27_40, w_carry_27_40;
math_adder_carry_save CSA_27_40(.i_a(w_pp_21_6), .i_b(w_pp_22_5), .i_c(w_pp_23_4), .ow_sum(w_sum_27_40), .ow_c(w_carry_27_40));
wire w_sum_27_38, w_carry_27_38;
math_adder_carry_save CSA_27_38(.i_a(w_pp_24_3), .i_b(w_pp_25_2), .i_c(w_pp_26_1), .ow_sum(w_sum_27_38), .ow_c(w_carry_27_38));
wire w_sum_27_36, w_carry_27_36;
math_adder_carry_save CSA_27_36(.i_a(w_pp_27_0), .i_b(w_carry_26_52), .i_c(w_carry_26_50), .ow_sum(w_sum_27_36), .ow_c(w_carry_27_36));
wire w_sum_27_34, w_carry_27_34;
math_adder_carry_save CSA_27_34(.i_a(w_carry_26_48), .i_b(w_carry_26_46), .i_c(w_carry_26_44), .ow_sum(w_sum_27_34), .ow_c(w_carry_27_34));
wire w_sum_27_32, w_carry_27_32;
math_adder_carry_save CSA_27_32(.i_a(w_carry_26_42), .i_b(w_carry_26_40), .i_c(w_carry_26_38), .ow_sum(w_sum_27_32), .ow_c(w_carry_27_32));
wire w_sum_27_30, w_carry_27_30;
math_adder_carry_save CSA_27_30(.i_a(w_carry_26_36), .i_b(w_carry_26_34), .i_c(w_carry_26_32), .ow_sum(w_sum_27_30), .ow_c(w_carry_27_30));
wire w_sum_27_28, w_carry_27_28;
math_adder_carry_save CSA_27_28(.i_a(w_carry_26_30), .i_b(w_carry_26_28), .i_c(w_carry_26_26), .ow_sum(w_sum_27_28), .ow_c(w_carry_27_28));
wire w_sum_27_26, w_carry_27_26;
math_adder_carry_save CSA_27_26(.i_a(w_carry_26_24), .i_b(w_carry_26_22), .i_c(w_carry_26_20), .ow_sum(w_sum_27_26), .ow_c(w_carry_27_26));
wire w_sum_27_24, w_carry_27_24;
math_adder_carry_save CSA_27_24(.i_a(w_carry_26_18), .i_b(w_carry_26_16), .i_c(w_carry_26_14), .ow_sum(w_sum_27_24), .ow_c(w_carry_27_24));
wire w_sum_27_22, w_carry_27_22;
math_adder_carry_save CSA_27_22(.i_a(w_carry_26_12), .i_b(w_carry_26_10), .i_c(w_carry_26_8), .ow_sum(w_sum_27_22), .ow_c(w_carry_27_22));
wire w_sum_27_20, w_carry_27_20;
math_adder_carry_save CSA_27_20(.i_a(w_carry_26_6), .i_b(w_carry_26_4), .i_c(w_carry_26_2), .ow_sum(w_sum_27_20), .ow_c(w_carry_27_20));
wire w_sum_27_18, w_carry_27_18;
math_adder_carry_save CSA_27_18(.i_a(w_sum_27_54), .i_b(w_sum_27_52), .i_c(w_sum_27_50), .ow_sum(w_sum_27_18), .ow_c(w_carry_27_18));
wire w_sum_27_16, w_carry_27_16;
math_adder_carry_save CSA_27_16(.i_a(w_sum_27_48), .i_b(w_sum_27_46), .i_c(w_sum_27_44), .ow_sum(w_sum_27_16), .ow_c(w_carry_27_16));
wire w_sum_27_14, w_carry_27_14;
math_adder_carry_save CSA_27_14(.i_a(w_sum_27_42), .i_b(w_sum_27_40), .i_c(w_sum_27_38), .ow_sum(w_sum_27_14), .ow_c(w_carry_27_14));
wire w_sum_27_12, w_carry_27_12;
math_adder_carry_save CSA_27_12(.i_a(w_sum_27_36), .i_b(w_sum_27_34), .i_c(w_sum_27_32), .ow_sum(w_sum_27_12), .ow_c(w_carry_27_12));
wire w_sum_27_10, w_carry_27_10;
math_adder_carry_save CSA_27_10(.i_a(w_sum_27_30), .i_b(w_sum_27_28), .i_c(w_sum_27_26), .ow_sum(w_sum_27_10), .ow_c(w_carry_27_10));
wire w_sum_27_8, w_carry_27_8;
math_adder_carry_save CSA_27_8(.i_a(w_sum_27_24), .i_b(w_sum_27_22), .i_c(w_sum_27_20), .ow_sum(w_sum_27_8), .ow_c(w_carry_27_8));
wire w_sum_27_6, w_carry_27_6;
math_adder_carry_save CSA_27_6(.i_a(w_sum_27_18), .i_b(w_sum_27_16), .i_c(w_sum_27_14), .ow_sum(w_sum_27_6), .ow_c(w_carry_27_6));
wire w_sum_27_4, w_carry_27_4;
math_adder_carry_save CSA_27_4(.i_a(w_sum_27_12), .i_b(w_sum_27_10), .i_c(w_sum_27_8), .ow_sum(w_sum_27_4), .ow_c(w_carry_27_4));
wire w_sum_27_2, w_carry_27_2;
math_adder_half HA_27_2(.i_a(w_sum_27_6), .i_b(w_sum_27_4), .ow_sum(w_sum_27_2), .ow_c(w_carry_27_2));
wire w_sum_28_56, w_carry_28_56;
math_adder_carry_save CSA_28_56(.i_a(w_pp_0_28), .i_b(w_pp_1_27), .i_c(w_pp_2_26), .ow_sum(w_sum_28_56), .ow_c(w_carry_28_56));
wire w_sum_28_54, w_carry_28_54;
math_adder_carry_save CSA_28_54(.i_a(w_pp_3_25), .i_b(w_pp_4_24), .i_c(w_pp_5_23), .ow_sum(w_sum_28_54), .ow_c(w_carry_28_54));
wire w_sum_28_52, w_carry_28_52;
math_adder_carry_save CSA_28_52(.i_a(w_pp_6_22), .i_b(w_pp_7_21), .i_c(w_pp_8_20), .ow_sum(w_sum_28_52), .ow_c(w_carry_28_52));
wire w_sum_28_50, w_carry_28_50;
math_adder_carry_save CSA_28_50(.i_a(w_pp_9_19), .i_b(w_pp_10_18), .i_c(w_pp_11_17), .ow_sum(w_sum_28_50), .ow_c(w_carry_28_50));
wire w_sum_28_48, w_carry_28_48;
math_adder_carry_save CSA_28_48(.i_a(w_pp_12_16), .i_b(w_pp_13_15), .i_c(w_pp_14_14), .ow_sum(w_sum_28_48), .ow_c(w_carry_28_48));
wire w_sum_28_46, w_carry_28_46;
math_adder_carry_save CSA_28_46(.i_a(w_pp_15_13), .i_b(w_pp_16_12), .i_c(w_pp_17_11), .ow_sum(w_sum_28_46), .ow_c(w_carry_28_46));
wire w_sum_28_44, w_carry_28_44;
math_adder_carry_save CSA_28_44(.i_a(w_pp_18_10), .i_b(w_pp_19_9), .i_c(w_pp_20_8), .ow_sum(w_sum_28_44), .ow_c(w_carry_28_44));
wire w_sum_28_42, w_carry_28_42;
math_adder_carry_save CSA_28_42(.i_a(w_pp_21_7), .i_b(w_pp_22_6), .i_c(w_pp_23_5), .ow_sum(w_sum_28_42), .ow_c(w_carry_28_42));
wire w_sum_28_40, w_carry_28_40;
math_adder_carry_save CSA_28_40(.i_a(w_pp_24_4), .i_b(w_pp_25_3), .i_c(w_pp_26_2), .ow_sum(w_sum_28_40), .ow_c(w_carry_28_40));
wire w_sum_28_38, w_carry_28_38;
math_adder_carry_save CSA_28_38(.i_a(w_pp_27_1), .i_b(w_pp_28_0), .i_c(w_carry_27_54), .ow_sum(w_sum_28_38), .ow_c(w_carry_28_38));
wire w_sum_28_36, w_carry_28_36;
math_adder_carry_save CSA_28_36(.i_a(w_carry_27_52), .i_b(w_carry_27_50), .i_c(w_carry_27_48), .ow_sum(w_sum_28_36), .ow_c(w_carry_28_36));
wire w_sum_28_34, w_carry_28_34;
math_adder_carry_save CSA_28_34(.i_a(w_carry_27_46), .i_b(w_carry_27_44), .i_c(w_carry_27_42), .ow_sum(w_sum_28_34), .ow_c(w_carry_28_34));
wire w_sum_28_32, w_carry_28_32;
math_adder_carry_save CSA_28_32(.i_a(w_carry_27_40), .i_b(w_carry_27_38), .i_c(w_carry_27_36), .ow_sum(w_sum_28_32), .ow_c(w_carry_28_32));
wire w_sum_28_30, w_carry_28_30;
math_adder_carry_save CSA_28_30(.i_a(w_carry_27_34), .i_b(w_carry_27_32), .i_c(w_carry_27_30), .ow_sum(w_sum_28_30), .ow_c(w_carry_28_30));
wire w_sum_28_28, w_carry_28_28;
math_adder_carry_save CSA_28_28(.i_a(w_carry_27_28), .i_b(w_carry_27_26), .i_c(w_carry_27_24), .ow_sum(w_sum_28_28), .ow_c(w_carry_28_28));
wire w_sum_28_26, w_carry_28_26;
math_adder_carry_save CSA_28_26(.i_a(w_carry_27_22), .i_b(w_carry_27_20), .i_c(w_carry_27_18), .ow_sum(w_sum_28_26), .ow_c(w_carry_28_26));
wire w_sum_28_24, w_carry_28_24;
math_adder_carry_save CSA_28_24(.i_a(w_carry_27_16), .i_b(w_carry_27_14), .i_c(w_carry_27_12), .ow_sum(w_sum_28_24), .ow_c(w_carry_28_24));
wire w_sum_28_22, w_carry_28_22;
math_adder_carry_save CSA_28_22(.i_a(w_carry_27_10), .i_b(w_carry_27_8), .i_c(w_carry_27_6), .ow_sum(w_sum_28_22), .ow_c(w_carry_28_22));
wire w_sum_28_20, w_carry_28_20;
math_adder_carry_save CSA_28_20(.i_a(w_carry_27_4), .i_b(w_carry_27_2), .i_c(w_sum_28_56), .ow_sum(w_sum_28_20), .ow_c(w_carry_28_20));
wire w_sum_28_18, w_carry_28_18;
math_adder_carry_save CSA_28_18(.i_a(w_sum_28_54), .i_b(w_sum_28_52), .i_c(w_sum_28_50), .ow_sum(w_sum_28_18), .ow_c(w_carry_28_18));
wire w_sum_28_16, w_carry_28_16;
math_adder_carry_save CSA_28_16(.i_a(w_sum_28_48), .i_b(w_sum_28_46), .i_c(w_sum_28_44), .ow_sum(w_sum_28_16), .ow_c(w_carry_28_16));
wire w_sum_28_14, w_carry_28_14;
math_adder_carry_save CSA_28_14(.i_a(w_sum_28_42), .i_b(w_sum_28_40), .i_c(w_sum_28_38), .ow_sum(w_sum_28_14), .ow_c(w_carry_28_14));
wire w_sum_28_12, w_carry_28_12;
math_adder_carry_save CSA_28_12(.i_a(w_sum_28_36), .i_b(w_sum_28_34), .i_c(w_sum_28_32), .ow_sum(w_sum_28_12), .ow_c(w_carry_28_12));
wire w_sum_28_10, w_carry_28_10;
math_adder_carry_save CSA_28_10(.i_a(w_sum_28_30), .i_b(w_sum_28_28), .i_c(w_sum_28_26), .ow_sum(w_sum_28_10), .ow_c(w_carry_28_10));
wire w_sum_28_8, w_carry_28_8;
math_adder_carry_save CSA_28_8(.i_a(w_sum_28_24), .i_b(w_sum_28_22), .i_c(w_sum_28_20), .ow_sum(w_sum_28_8), .ow_c(w_carry_28_8));
wire w_sum_28_6, w_carry_28_6;
math_adder_carry_save CSA_28_6(.i_a(w_sum_28_18), .i_b(w_sum_28_16), .i_c(w_sum_28_14), .ow_sum(w_sum_28_6), .ow_c(w_carry_28_6));
wire w_sum_28_4, w_carry_28_4;
math_adder_carry_save CSA_28_4(.i_a(w_sum_28_12), .i_b(w_sum_28_10), .i_c(w_sum_28_8), .ow_sum(w_sum_28_4), .ow_c(w_carry_28_4));
wire w_sum_28_2, w_carry_28_2;
math_adder_half HA_28_2(.i_a(w_sum_28_6), .i_b(w_sum_28_4), .ow_sum(w_sum_28_2), .ow_c(w_carry_28_2));
wire w_sum_29_58, w_carry_29_58;
math_adder_carry_save CSA_29_58(.i_a(w_pp_0_29), .i_b(w_pp_1_28), .i_c(w_pp_2_27), .ow_sum(w_sum_29_58), .ow_c(w_carry_29_58));
wire w_sum_29_56, w_carry_29_56;
math_adder_carry_save CSA_29_56(.i_a(w_pp_3_26), .i_b(w_pp_4_25), .i_c(w_pp_5_24), .ow_sum(w_sum_29_56), .ow_c(w_carry_29_56));
wire w_sum_29_54, w_carry_29_54;
math_adder_carry_save CSA_29_54(.i_a(w_pp_6_23), .i_b(w_pp_7_22), .i_c(w_pp_8_21), .ow_sum(w_sum_29_54), .ow_c(w_carry_29_54));
wire w_sum_29_52, w_carry_29_52;
math_adder_carry_save CSA_29_52(.i_a(w_pp_9_20), .i_b(w_pp_10_19), .i_c(w_pp_11_18), .ow_sum(w_sum_29_52), .ow_c(w_carry_29_52));
wire w_sum_29_50, w_carry_29_50;
math_adder_carry_save CSA_29_50(.i_a(w_pp_12_17), .i_b(w_pp_13_16), .i_c(w_pp_14_15), .ow_sum(w_sum_29_50), .ow_c(w_carry_29_50));
wire w_sum_29_48, w_carry_29_48;
math_adder_carry_save CSA_29_48(.i_a(w_pp_15_14), .i_b(w_pp_16_13), .i_c(w_pp_17_12), .ow_sum(w_sum_29_48), .ow_c(w_carry_29_48));
wire w_sum_29_46, w_carry_29_46;
math_adder_carry_save CSA_29_46(.i_a(w_pp_18_11), .i_b(w_pp_19_10), .i_c(w_pp_20_9), .ow_sum(w_sum_29_46), .ow_c(w_carry_29_46));
wire w_sum_29_44, w_carry_29_44;
math_adder_carry_save CSA_29_44(.i_a(w_pp_21_8), .i_b(w_pp_22_7), .i_c(w_pp_23_6), .ow_sum(w_sum_29_44), .ow_c(w_carry_29_44));
wire w_sum_29_42, w_carry_29_42;
math_adder_carry_save CSA_29_42(.i_a(w_pp_24_5), .i_b(w_pp_25_4), .i_c(w_pp_26_3), .ow_sum(w_sum_29_42), .ow_c(w_carry_29_42));
wire w_sum_29_40, w_carry_29_40;
math_adder_carry_save CSA_29_40(.i_a(w_pp_27_2), .i_b(w_pp_28_1), .i_c(w_pp_29_0), .ow_sum(w_sum_29_40), .ow_c(w_carry_29_40));
wire w_sum_29_38, w_carry_29_38;
math_adder_carry_save CSA_29_38(.i_a(w_carry_28_56), .i_b(w_carry_28_54), .i_c(w_carry_28_52), .ow_sum(w_sum_29_38), .ow_c(w_carry_29_38));
wire w_sum_29_36, w_carry_29_36;
math_adder_carry_save CSA_29_36(.i_a(w_carry_28_50), .i_b(w_carry_28_48), .i_c(w_carry_28_46), .ow_sum(w_sum_29_36), .ow_c(w_carry_29_36));
wire w_sum_29_34, w_carry_29_34;
math_adder_carry_save CSA_29_34(.i_a(w_carry_28_44), .i_b(w_carry_28_42), .i_c(w_carry_28_40), .ow_sum(w_sum_29_34), .ow_c(w_carry_29_34));
wire w_sum_29_32, w_carry_29_32;
math_adder_carry_save CSA_29_32(.i_a(w_carry_28_38), .i_b(w_carry_28_36), .i_c(w_carry_28_34), .ow_sum(w_sum_29_32), .ow_c(w_carry_29_32));
wire w_sum_29_30, w_carry_29_30;
math_adder_carry_save CSA_29_30(.i_a(w_carry_28_32), .i_b(w_carry_28_30), .i_c(w_carry_28_28), .ow_sum(w_sum_29_30), .ow_c(w_carry_29_30));
wire w_sum_29_28, w_carry_29_28;
math_adder_carry_save CSA_29_28(.i_a(w_carry_28_26), .i_b(w_carry_28_24), .i_c(w_carry_28_22), .ow_sum(w_sum_29_28), .ow_c(w_carry_29_28));
wire w_sum_29_26, w_carry_29_26;
math_adder_carry_save CSA_29_26(.i_a(w_carry_28_20), .i_b(w_carry_28_18), .i_c(w_carry_28_16), .ow_sum(w_sum_29_26), .ow_c(w_carry_29_26));
wire w_sum_29_24, w_carry_29_24;
math_adder_carry_save CSA_29_24(.i_a(w_carry_28_14), .i_b(w_carry_28_12), .i_c(w_carry_28_10), .ow_sum(w_sum_29_24), .ow_c(w_carry_29_24));
wire w_sum_29_22, w_carry_29_22;
math_adder_carry_save CSA_29_22(.i_a(w_carry_28_8), .i_b(w_carry_28_6), .i_c(w_carry_28_4), .ow_sum(w_sum_29_22), .ow_c(w_carry_29_22));
wire w_sum_29_20, w_carry_29_20;
math_adder_carry_save CSA_29_20(.i_a(w_carry_28_2), .i_b(w_sum_29_58), .i_c(w_sum_29_56), .ow_sum(w_sum_29_20), .ow_c(w_carry_29_20));
wire w_sum_29_18, w_carry_29_18;
math_adder_carry_save CSA_29_18(.i_a(w_sum_29_54), .i_b(w_sum_29_52), .i_c(w_sum_29_50), .ow_sum(w_sum_29_18), .ow_c(w_carry_29_18));
wire w_sum_29_16, w_carry_29_16;
math_adder_carry_save CSA_29_16(.i_a(w_sum_29_48), .i_b(w_sum_29_46), .i_c(w_sum_29_44), .ow_sum(w_sum_29_16), .ow_c(w_carry_29_16));
wire w_sum_29_14, w_carry_29_14;
math_adder_carry_save CSA_29_14(.i_a(w_sum_29_42), .i_b(w_sum_29_40), .i_c(w_sum_29_38), .ow_sum(w_sum_29_14), .ow_c(w_carry_29_14));
wire w_sum_29_12, w_carry_29_12;
math_adder_carry_save CSA_29_12(.i_a(w_sum_29_36), .i_b(w_sum_29_34), .i_c(w_sum_29_32), .ow_sum(w_sum_29_12), .ow_c(w_carry_29_12));
wire w_sum_29_10, w_carry_29_10;
math_adder_carry_save CSA_29_10(.i_a(w_sum_29_30), .i_b(w_sum_29_28), .i_c(w_sum_29_26), .ow_sum(w_sum_29_10), .ow_c(w_carry_29_10));
wire w_sum_29_8, w_carry_29_8;
math_adder_carry_save CSA_29_8(.i_a(w_sum_29_24), .i_b(w_sum_29_22), .i_c(w_sum_29_20), .ow_sum(w_sum_29_8), .ow_c(w_carry_29_8));
wire w_sum_29_6, w_carry_29_6;
math_adder_carry_save CSA_29_6(.i_a(w_sum_29_18), .i_b(w_sum_29_16), .i_c(w_sum_29_14), .ow_sum(w_sum_29_6), .ow_c(w_carry_29_6));
wire w_sum_29_4, w_carry_29_4;
math_adder_carry_save CSA_29_4(.i_a(w_sum_29_12), .i_b(w_sum_29_10), .i_c(w_sum_29_8), .ow_sum(w_sum_29_4), .ow_c(w_carry_29_4));
wire w_sum_29_2, w_carry_29_2;
math_adder_half HA_29_2(.i_a(w_sum_29_6), .i_b(w_sum_29_4), .ow_sum(w_sum_29_2), .ow_c(w_carry_29_2));
wire w_sum_30_60, w_carry_30_60;
math_adder_carry_save CSA_30_60(.i_a(w_pp_0_30), .i_b(w_pp_1_29), .i_c(w_pp_2_28), .ow_sum(w_sum_30_60), .ow_c(w_carry_30_60));
wire w_sum_30_58, w_carry_30_58;
math_adder_carry_save CSA_30_58(.i_a(w_pp_3_27), .i_b(w_pp_4_26), .i_c(w_pp_5_25), .ow_sum(w_sum_30_58), .ow_c(w_carry_30_58));
wire w_sum_30_56, w_carry_30_56;
math_adder_carry_save CSA_30_56(.i_a(w_pp_6_24), .i_b(w_pp_7_23), .i_c(w_pp_8_22), .ow_sum(w_sum_30_56), .ow_c(w_carry_30_56));
wire w_sum_30_54, w_carry_30_54;
math_adder_carry_save CSA_30_54(.i_a(w_pp_9_21), .i_b(w_pp_10_20), .i_c(w_pp_11_19), .ow_sum(w_sum_30_54), .ow_c(w_carry_30_54));
wire w_sum_30_52, w_carry_30_52;
math_adder_carry_save CSA_30_52(.i_a(w_pp_12_18), .i_b(w_pp_13_17), .i_c(w_pp_14_16), .ow_sum(w_sum_30_52), .ow_c(w_carry_30_52));
wire w_sum_30_50, w_carry_30_50;
math_adder_carry_save CSA_30_50(.i_a(w_pp_15_15), .i_b(w_pp_16_14), .i_c(w_pp_17_13), .ow_sum(w_sum_30_50), .ow_c(w_carry_30_50));
wire w_sum_30_48, w_carry_30_48;
math_adder_carry_save CSA_30_48(.i_a(w_pp_18_12), .i_b(w_pp_19_11), .i_c(w_pp_20_10), .ow_sum(w_sum_30_48), .ow_c(w_carry_30_48));
wire w_sum_30_46, w_carry_30_46;
math_adder_carry_save CSA_30_46(.i_a(w_pp_21_9), .i_b(w_pp_22_8), .i_c(w_pp_23_7), .ow_sum(w_sum_30_46), .ow_c(w_carry_30_46));
wire w_sum_30_44, w_carry_30_44;
math_adder_carry_save CSA_30_44(.i_a(w_pp_24_6), .i_b(w_pp_25_5), .i_c(w_pp_26_4), .ow_sum(w_sum_30_44), .ow_c(w_carry_30_44));
wire w_sum_30_42, w_carry_30_42;
math_adder_carry_save CSA_30_42(.i_a(w_pp_27_3), .i_b(w_pp_28_2), .i_c(w_pp_29_1), .ow_sum(w_sum_30_42), .ow_c(w_carry_30_42));
wire w_sum_30_40, w_carry_30_40;
math_adder_carry_save CSA_30_40(.i_a(w_pp_30_0), .i_b(w_carry_29_58), .i_c(w_carry_29_56), .ow_sum(w_sum_30_40), .ow_c(w_carry_30_40));
wire w_sum_30_38, w_carry_30_38;
math_adder_carry_save CSA_30_38(.i_a(w_carry_29_54), .i_b(w_carry_29_52), .i_c(w_carry_29_50), .ow_sum(w_sum_30_38), .ow_c(w_carry_30_38));
wire w_sum_30_36, w_carry_30_36;
math_adder_carry_save CSA_30_36(.i_a(w_carry_29_48), .i_b(w_carry_29_46), .i_c(w_carry_29_44), .ow_sum(w_sum_30_36), .ow_c(w_carry_30_36));
wire w_sum_30_34, w_carry_30_34;
math_adder_carry_save CSA_30_34(.i_a(w_carry_29_42), .i_b(w_carry_29_40), .i_c(w_carry_29_38), .ow_sum(w_sum_30_34), .ow_c(w_carry_30_34));
wire w_sum_30_32, w_carry_30_32;
math_adder_carry_save CSA_30_32(.i_a(w_carry_29_36), .i_b(w_carry_29_34), .i_c(w_carry_29_32), .ow_sum(w_sum_30_32), .ow_c(w_carry_30_32));
wire w_sum_30_30, w_carry_30_30;
math_adder_carry_save CSA_30_30(.i_a(w_carry_29_30), .i_b(w_carry_29_28), .i_c(w_carry_29_26), .ow_sum(w_sum_30_30), .ow_c(w_carry_30_30));
wire w_sum_30_28, w_carry_30_28;
math_adder_carry_save CSA_30_28(.i_a(w_carry_29_24), .i_b(w_carry_29_22), .i_c(w_carry_29_20), .ow_sum(w_sum_30_28), .ow_c(w_carry_30_28));
wire w_sum_30_26, w_carry_30_26;
math_adder_carry_save CSA_30_26(.i_a(w_carry_29_18), .i_b(w_carry_29_16), .i_c(w_carry_29_14), .ow_sum(w_sum_30_26), .ow_c(w_carry_30_26));
wire w_sum_30_24, w_carry_30_24;
math_adder_carry_save CSA_30_24(.i_a(w_carry_29_12), .i_b(w_carry_29_10), .i_c(w_carry_29_8), .ow_sum(w_sum_30_24), .ow_c(w_carry_30_24));
wire w_sum_30_22, w_carry_30_22;
math_adder_carry_save CSA_30_22(.i_a(w_carry_29_6), .i_b(w_carry_29_4), .i_c(w_carry_29_2), .ow_sum(w_sum_30_22), .ow_c(w_carry_30_22));
wire w_sum_30_20, w_carry_30_20;
math_adder_carry_save CSA_30_20(.i_a(w_sum_30_60), .i_b(w_sum_30_58), .i_c(w_sum_30_56), .ow_sum(w_sum_30_20), .ow_c(w_carry_30_20));
wire w_sum_30_18, w_carry_30_18;
math_adder_carry_save CSA_30_18(.i_a(w_sum_30_54), .i_b(w_sum_30_52), .i_c(w_sum_30_50), .ow_sum(w_sum_30_18), .ow_c(w_carry_30_18));
wire w_sum_30_16, w_carry_30_16;
math_adder_carry_save CSA_30_16(.i_a(w_sum_30_48), .i_b(w_sum_30_46), .i_c(w_sum_30_44), .ow_sum(w_sum_30_16), .ow_c(w_carry_30_16));
wire w_sum_30_14, w_carry_30_14;
math_adder_carry_save CSA_30_14(.i_a(w_sum_30_42), .i_b(w_sum_30_40), .i_c(w_sum_30_38), .ow_sum(w_sum_30_14), .ow_c(w_carry_30_14));
wire w_sum_30_12, w_carry_30_12;
math_adder_carry_save CSA_30_12(.i_a(w_sum_30_36), .i_b(w_sum_30_34), .i_c(w_sum_30_32), .ow_sum(w_sum_30_12), .ow_c(w_carry_30_12));
wire w_sum_30_10, w_carry_30_10;
math_adder_carry_save CSA_30_10(.i_a(w_sum_30_30), .i_b(w_sum_30_28), .i_c(w_sum_30_26), .ow_sum(w_sum_30_10), .ow_c(w_carry_30_10));
wire w_sum_30_8, w_carry_30_8;
math_adder_carry_save CSA_30_8(.i_a(w_sum_30_24), .i_b(w_sum_30_22), .i_c(w_sum_30_20), .ow_sum(w_sum_30_8), .ow_c(w_carry_30_8));
wire w_sum_30_6, w_carry_30_6;
math_adder_carry_save CSA_30_6(.i_a(w_sum_30_18), .i_b(w_sum_30_16), .i_c(w_sum_30_14), .ow_sum(w_sum_30_6), .ow_c(w_carry_30_6));
wire w_sum_30_4, w_carry_30_4;
math_adder_carry_save CSA_30_4(.i_a(w_sum_30_12), .i_b(w_sum_30_10), .i_c(w_sum_30_8), .ow_sum(w_sum_30_4), .ow_c(w_carry_30_4));
wire w_sum_30_2, w_carry_30_2;
math_adder_half HA_30_2(.i_a(w_sum_30_6), .i_b(w_sum_30_4), .ow_sum(w_sum_30_2), .ow_c(w_carry_30_2));
wire w_sum_31_62, w_carry_31_62;
math_adder_carry_save CSA_31_62(.i_a(w_pp_0_31), .i_b(w_pp_1_30), .i_c(w_pp_2_29), .ow_sum(w_sum_31_62), .ow_c(w_carry_31_62));
wire w_sum_31_60, w_carry_31_60;
math_adder_carry_save CSA_31_60(.i_a(w_pp_3_28), .i_b(w_pp_4_27), .i_c(w_pp_5_26), .ow_sum(w_sum_31_60), .ow_c(w_carry_31_60));
wire w_sum_31_58, w_carry_31_58;
math_adder_carry_save CSA_31_58(.i_a(w_pp_6_25), .i_b(w_pp_7_24), .i_c(w_pp_8_23), .ow_sum(w_sum_31_58), .ow_c(w_carry_31_58));
wire w_sum_31_56, w_carry_31_56;
math_adder_carry_save CSA_31_56(.i_a(w_pp_9_22), .i_b(w_pp_10_21), .i_c(w_pp_11_20), .ow_sum(w_sum_31_56), .ow_c(w_carry_31_56));
wire w_sum_31_54, w_carry_31_54;
math_adder_carry_save CSA_31_54(.i_a(w_pp_12_19), .i_b(w_pp_13_18), .i_c(w_pp_14_17), .ow_sum(w_sum_31_54), .ow_c(w_carry_31_54));
wire w_sum_31_52, w_carry_31_52;
math_adder_carry_save CSA_31_52(.i_a(w_pp_15_16), .i_b(w_pp_16_15), .i_c(w_pp_17_14), .ow_sum(w_sum_31_52), .ow_c(w_carry_31_52));
wire w_sum_31_50, w_carry_31_50;
math_adder_carry_save CSA_31_50(.i_a(w_pp_18_13), .i_b(w_pp_19_12), .i_c(w_pp_20_11), .ow_sum(w_sum_31_50), .ow_c(w_carry_31_50));
wire w_sum_31_48, w_carry_31_48;
math_adder_carry_save CSA_31_48(.i_a(w_pp_21_10), .i_b(w_pp_22_9), .i_c(w_pp_23_8), .ow_sum(w_sum_31_48), .ow_c(w_carry_31_48));
wire w_sum_31_46, w_carry_31_46;
math_adder_carry_save CSA_31_46(.i_a(w_pp_24_7), .i_b(w_pp_25_6), .i_c(w_pp_26_5), .ow_sum(w_sum_31_46), .ow_c(w_carry_31_46));
wire w_sum_31_44, w_carry_31_44;
math_adder_carry_save CSA_31_44(.i_a(w_pp_27_4), .i_b(w_pp_28_3), .i_c(w_pp_29_2), .ow_sum(w_sum_31_44), .ow_c(w_carry_31_44));
wire w_sum_31_42, w_carry_31_42;
math_adder_carry_save CSA_31_42(.i_a(w_pp_30_1), .i_b(w_pp_31_0), .i_c(w_carry_30_60), .ow_sum(w_sum_31_42), .ow_c(w_carry_31_42));
wire w_sum_31_40, w_carry_31_40;
math_adder_carry_save CSA_31_40(.i_a(w_carry_30_58), .i_b(w_carry_30_56), .i_c(w_carry_30_54), .ow_sum(w_sum_31_40), .ow_c(w_carry_31_40));
wire w_sum_31_38, w_carry_31_38;
math_adder_carry_save CSA_31_38(.i_a(w_carry_30_52), .i_b(w_carry_30_50), .i_c(w_carry_30_48), .ow_sum(w_sum_31_38), .ow_c(w_carry_31_38));
wire w_sum_31_36, w_carry_31_36;
math_adder_carry_save CSA_31_36(.i_a(w_carry_30_46), .i_b(w_carry_30_44), .i_c(w_carry_30_42), .ow_sum(w_sum_31_36), .ow_c(w_carry_31_36));
wire w_sum_31_34, w_carry_31_34;
math_adder_carry_save CSA_31_34(.i_a(w_carry_30_40), .i_b(w_carry_30_38), .i_c(w_carry_30_36), .ow_sum(w_sum_31_34), .ow_c(w_carry_31_34));
wire w_sum_31_32, w_carry_31_32;
math_adder_carry_save CSA_31_32(.i_a(w_carry_30_34), .i_b(w_carry_30_32), .i_c(w_carry_30_30), .ow_sum(w_sum_31_32), .ow_c(w_carry_31_32));
wire w_sum_31_30, w_carry_31_30;
math_adder_carry_save CSA_31_30(.i_a(w_carry_30_28), .i_b(w_carry_30_26), .i_c(w_carry_30_24), .ow_sum(w_sum_31_30), .ow_c(w_carry_31_30));
wire w_sum_31_28, w_carry_31_28;
math_adder_carry_save CSA_31_28(.i_a(w_carry_30_22), .i_b(w_carry_30_20), .i_c(w_carry_30_18), .ow_sum(w_sum_31_28), .ow_c(w_carry_31_28));
wire w_sum_31_26, w_carry_31_26;
math_adder_carry_save CSA_31_26(.i_a(w_carry_30_16), .i_b(w_carry_30_14), .i_c(w_carry_30_12), .ow_sum(w_sum_31_26), .ow_c(w_carry_31_26));
wire w_sum_31_24, w_carry_31_24;
math_adder_carry_save CSA_31_24(.i_a(w_carry_30_10), .i_b(w_carry_30_8), .i_c(w_carry_30_6), .ow_sum(w_sum_31_24), .ow_c(w_carry_31_24));
wire w_sum_31_22, w_carry_31_22;
math_adder_carry_save CSA_31_22(.i_a(w_carry_30_4), .i_b(w_carry_30_2), .i_c(w_sum_31_62), .ow_sum(w_sum_31_22), .ow_c(w_carry_31_22));
wire w_sum_31_20, w_carry_31_20;
math_adder_carry_save CSA_31_20(.i_a(w_sum_31_60), .i_b(w_sum_31_58), .i_c(w_sum_31_56), .ow_sum(w_sum_31_20), .ow_c(w_carry_31_20));
wire w_sum_31_18, w_carry_31_18;
math_adder_carry_save CSA_31_18(.i_a(w_sum_31_54), .i_b(w_sum_31_52), .i_c(w_sum_31_50), .ow_sum(w_sum_31_18), .ow_c(w_carry_31_18));
wire w_sum_31_16, w_carry_31_16;
math_adder_carry_save CSA_31_16(.i_a(w_sum_31_48), .i_b(w_sum_31_46), .i_c(w_sum_31_44), .ow_sum(w_sum_31_16), .ow_c(w_carry_31_16));
wire w_sum_31_14, w_carry_31_14;
math_adder_carry_save CSA_31_14(.i_a(w_sum_31_42), .i_b(w_sum_31_40), .i_c(w_sum_31_38), .ow_sum(w_sum_31_14), .ow_c(w_carry_31_14));
wire w_sum_31_12, w_carry_31_12;
math_adder_carry_save CSA_31_12(.i_a(w_sum_31_36), .i_b(w_sum_31_34), .i_c(w_sum_31_32), .ow_sum(w_sum_31_12), .ow_c(w_carry_31_12));
wire w_sum_31_10, w_carry_31_10;
math_adder_carry_save CSA_31_10(.i_a(w_sum_31_30), .i_b(w_sum_31_28), .i_c(w_sum_31_26), .ow_sum(w_sum_31_10), .ow_c(w_carry_31_10));
wire w_sum_31_8, w_carry_31_8;
math_adder_carry_save CSA_31_8(.i_a(w_sum_31_24), .i_b(w_sum_31_22), .i_c(w_sum_31_20), .ow_sum(w_sum_31_8), .ow_c(w_carry_31_8));
wire w_sum_31_6, w_carry_31_6;
math_adder_carry_save CSA_31_6(.i_a(w_sum_31_18), .i_b(w_sum_31_16), .i_c(w_sum_31_14), .ow_sum(w_sum_31_6), .ow_c(w_carry_31_6));
wire w_sum_31_4, w_carry_31_4;
math_adder_carry_save CSA_31_4(.i_a(w_sum_31_12), .i_b(w_sum_31_10), .i_c(w_sum_31_8), .ow_sum(w_sum_31_4), .ow_c(w_carry_31_4));
wire w_sum_31_2, w_carry_31_2;
math_adder_half HA_31_2(.i_a(w_sum_31_6), .i_b(w_sum_31_4), .ow_sum(w_sum_31_2), .ow_c(w_carry_31_2));
wire w_sum_32_62, w_carry_32_62;
math_adder_carry_save CSA_32_62(.i_a(w_pp_1_31), .i_b(w_pp_2_30), .i_c(w_pp_3_29), .ow_sum(w_sum_32_62), .ow_c(w_carry_32_62));
wire w_sum_32_60, w_carry_32_60;
math_adder_carry_save CSA_32_60(.i_a(w_pp_4_28), .i_b(w_pp_5_27), .i_c(w_pp_6_26), .ow_sum(w_sum_32_60), .ow_c(w_carry_32_60));
wire w_sum_32_58, w_carry_32_58;
math_adder_carry_save CSA_32_58(.i_a(w_pp_7_25), .i_b(w_pp_8_24), .i_c(w_pp_9_23), .ow_sum(w_sum_32_58), .ow_c(w_carry_32_58));
wire w_sum_32_56, w_carry_32_56;
math_adder_carry_save CSA_32_56(.i_a(w_pp_10_22), .i_b(w_pp_11_21), .i_c(w_pp_12_20), .ow_sum(w_sum_32_56), .ow_c(w_carry_32_56));
wire w_sum_32_54, w_carry_32_54;
math_adder_carry_save CSA_32_54(.i_a(w_pp_13_19), .i_b(w_pp_14_18), .i_c(w_pp_15_17), .ow_sum(w_sum_32_54), .ow_c(w_carry_32_54));
wire w_sum_32_52, w_carry_32_52;
math_adder_carry_save CSA_32_52(.i_a(w_pp_16_16), .i_b(w_pp_17_15), .i_c(w_pp_18_14), .ow_sum(w_sum_32_52), .ow_c(w_carry_32_52));
wire w_sum_32_50, w_carry_32_50;
math_adder_carry_save CSA_32_50(.i_a(w_pp_19_13), .i_b(w_pp_20_12), .i_c(w_pp_21_11), .ow_sum(w_sum_32_50), .ow_c(w_carry_32_50));
wire w_sum_32_48, w_carry_32_48;
math_adder_carry_save CSA_32_48(.i_a(w_pp_22_10), .i_b(w_pp_23_9), .i_c(w_pp_24_8), .ow_sum(w_sum_32_48), .ow_c(w_carry_32_48));
wire w_sum_32_46, w_carry_32_46;
math_adder_carry_save CSA_32_46(.i_a(w_pp_25_7), .i_b(w_pp_26_6), .i_c(w_pp_27_5), .ow_sum(w_sum_32_46), .ow_c(w_carry_32_46));
wire w_sum_32_44, w_carry_32_44;
math_adder_carry_save CSA_32_44(.i_a(w_pp_28_4), .i_b(w_pp_29_3), .i_c(w_pp_30_2), .ow_sum(w_sum_32_44), .ow_c(w_carry_32_44));
wire w_sum_32_42, w_carry_32_42;
math_adder_carry_save CSA_32_42(.i_a(w_pp_31_1), .i_b(w_carry_31_62), .i_c(w_carry_31_60), .ow_sum(w_sum_32_42), .ow_c(w_carry_32_42));
wire w_sum_32_40, w_carry_32_40;
math_adder_carry_save CSA_32_40(.i_a(w_carry_31_58), .i_b(w_carry_31_56), .i_c(w_carry_31_54), .ow_sum(w_sum_32_40), .ow_c(w_carry_32_40));
wire w_sum_32_38, w_carry_32_38;
math_adder_carry_save CSA_32_38(.i_a(w_carry_31_52), .i_b(w_carry_31_50), .i_c(w_carry_31_48), .ow_sum(w_sum_32_38), .ow_c(w_carry_32_38));
wire w_sum_32_36, w_carry_32_36;
math_adder_carry_save CSA_32_36(.i_a(w_carry_31_46), .i_b(w_carry_31_44), .i_c(w_carry_31_42), .ow_sum(w_sum_32_36), .ow_c(w_carry_32_36));
wire w_sum_32_34, w_carry_32_34;
math_adder_carry_save CSA_32_34(.i_a(w_carry_31_40), .i_b(w_carry_31_38), .i_c(w_carry_31_36), .ow_sum(w_sum_32_34), .ow_c(w_carry_32_34));
wire w_sum_32_32, w_carry_32_32;
math_adder_carry_save CSA_32_32(.i_a(w_carry_31_34), .i_b(w_carry_31_32), .i_c(w_carry_31_30), .ow_sum(w_sum_32_32), .ow_c(w_carry_32_32));
wire w_sum_32_30, w_carry_32_30;
math_adder_carry_save CSA_32_30(.i_a(w_carry_31_28), .i_b(w_carry_31_26), .i_c(w_carry_31_24), .ow_sum(w_sum_32_30), .ow_c(w_carry_32_30));
wire w_sum_32_28, w_carry_32_28;
math_adder_carry_save CSA_32_28(.i_a(w_carry_31_22), .i_b(w_carry_31_20), .i_c(w_carry_31_18), .ow_sum(w_sum_32_28), .ow_c(w_carry_32_28));
wire w_sum_32_26, w_carry_32_26;
math_adder_carry_save CSA_32_26(.i_a(w_carry_31_16), .i_b(w_carry_31_14), .i_c(w_carry_31_12), .ow_sum(w_sum_32_26), .ow_c(w_carry_32_26));
wire w_sum_32_24, w_carry_32_24;
math_adder_carry_save CSA_32_24(.i_a(w_carry_31_10), .i_b(w_carry_31_8), .i_c(w_carry_31_6), .ow_sum(w_sum_32_24), .ow_c(w_carry_32_24));
wire w_sum_32_22, w_carry_32_22;
math_adder_carry_save CSA_32_22(.i_a(w_carry_31_4), .i_b(w_carry_31_2), .i_c(w_sum_32_62), .ow_sum(w_sum_32_22), .ow_c(w_carry_32_22));
wire w_sum_32_20, w_carry_32_20;
math_adder_carry_save CSA_32_20(.i_a(w_sum_32_60), .i_b(w_sum_32_58), .i_c(w_sum_32_56), .ow_sum(w_sum_32_20), .ow_c(w_carry_32_20));
wire w_sum_32_18, w_carry_32_18;
math_adder_carry_save CSA_32_18(.i_a(w_sum_32_54), .i_b(w_sum_32_52), .i_c(w_sum_32_50), .ow_sum(w_sum_32_18), .ow_c(w_carry_32_18));
wire w_sum_32_16, w_carry_32_16;
math_adder_carry_save CSA_32_16(.i_a(w_sum_32_48), .i_b(w_sum_32_46), .i_c(w_sum_32_44), .ow_sum(w_sum_32_16), .ow_c(w_carry_32_16));
wire w_sum_32_14, w_carry_32_14;
math_adder_carry_save CSA_32_14(.i_a(w_sum_32_42), .i_b(w_sum_32_40), .i_c(w_sum_32_38), .ow_sum(w_sum_32_14), .ow_c(w_carry_32_14));
wire w_sum_32_12, w_carry_32_12;
math_adder_carry_save CSA_32_12(.i_a(w_sum_32_36), .i_b(w_sum_32_34), .i_c(w_sum_32_32), .ow_sum(w_sum_32_12), .ow_c(w_carry_32_12));
wire w_sum_32_10, w_carry_32_10;
math_adder_carry_save CSA_32_10(.i_a(w_sum_32_30), .i_b(w_sum_32_28), .i_c(w_sum_32_26), .ow_sum(w_sum_32_10), .ow_c(w_carry_32_10));
wire w_sum_32_8, w_carry_32_8;
math_adder_carry_save CSA_32_8(.i_a(w_sum_32_24), .i_b(w_sum_32_22), .i_c(w_sum_32_20), .ow_sum(w_sum_32_8), .ow_c(w_carry_32_8));
wire w_sum_32_6, w_carry_32_6;
math_adder_carry_save CSA_32_6(.i_a(w_sum_32_18), .i_b(w_sum_32_16), .i_c(w_sum_32_14), .ow_sum(w_sum_32_6), .ow_c(w_carry_32_6));
wire w_sum_32_4, w_carry_32_4;
math_adder_carry_save CSA_32_4(.i_a(w_sum_32_12), .i_b(w_sum_32_10), .i_c(w_sum_32_8), .ow_sum(w_sum_32_4), .ow_c(w_carry_32_4));
wire w_sum_32_2, w_carry_32_2;
math_adder_half HA_32_2(.i_a(w_sum_32_6), .i_b(w_sum_32_4), .ow_sum(w_sum_32_2), .ow_c(w_carry_32_2));
wire w_sum_33_61, w_carry_33_61;
math_adder_carry_save CSA_33_61(.i_a(w_pp_2_31), .i_b(w_pp_3_30), .i_c(w_pp_4_29), .ow_sum(w_sum_33_61), .ow_c(w_carry_33_61));
wire w_sum_33_59, w_carry_33_59;
math_adder_carry_save CSA_33_59(.i_a(w_pp_5_28), .i_b(w_pp_6_27), .i_c(w_pp_7_26), .ow_sum(w_sum_33_59), .ow_c(w_carry_33_59));
wire w_sum_33_57, w_carry_33_57;
math_adder_carry_save CSA_33_57(.i_a(w_pp_8_25), .i_b(w_pp_9_24), .i_c(w_pp_10_23), .ow_sum(w_sum_33_57), .ow_c(w_carry_33_57));
wire w_sum_33_55, w_carry_33_55;
math_adder_carry_save CSA_33_55(.i_a(w_pp_11_22), .i_b(w_pp_12_21), .i_c(w_pp_13_20), .ow_sum(w_sum_33_55), .ow_c(w_carry_33_55));
wire w_sum_33_53, w_carry_33_53;
math_adder_carry_save CSA_33_53(.i_a(w_pp_14_19), .i_b(w_pp_15_18), .i_c(w_pp_16_17), .ow_sum(w_sum_33_53), .ow_c(w_carry_33_53));
wire w_sum_33_51, w_carry_33_51;
math_adder_carry_save CSA_33_51(.i_a(w_pp_17_16), .i_b(w_pp_18_15), .i_c(w_pp_19_14), .ow_sum(w_sum_33_51), .ow_c(w_carry_33_51));
wire w_sum_33_49, w_carry_33_49;
math_adder_carry_save CSA_33_49(.i_a(w_pp_20_13), .i_b(w_pp_21_12), .i_c(w_pp_22_11), .ow_sum(w_sum_33_49), .ow_c(w_carry_33_49));
wire w_sum_33_47, w_carry_33_47;
math_adder_carry_save CSA_33_47(.i_a(w_pp_23_10), .i_b(w_pp_24_9), .i_c(w_pp_25_8), .ow_sum(w_sum_33_47), .ow_c(w_carry_33_47));
wire w_sum_33_45, w_carry_33_45;
math_adder_carry_save CSA_33_45(.i_a(w_pp_26_7), .i_b(w_pp_27_6), .i_c(w_pp_28_5), .ow_sum(w_sum_33_45), .ow_c(w_carry_33_45));
wire w_sum_33_43, w_carry_33_43;
math_adder_carry_save CSA_33_43(.i_a(w_pp_29_4), .i_b(w_pp_30_3), .i_c(w_pp_31_2), .ow_sum(w_sum_33_43), .ow_c(w_carry_33_43));
wire w_sum_33_41, w_carry_33_41;
math_adder_carry_save CSA_33_41(.i_a(w_carry_32_62), .i_b(w_carry_32_60), .i_c(w_carry_32_58), .ow_sum(w_sum_33_41), .ow_c(w_carry_33_41));
wire w_sum_33_39, w_carry_33_39;
math_adder_carry_save CSA_33_39(.i_a(w_carry_32_56), .i_b(w_carry_32_54), .i_c(w_carry_32_52), .ow_sum(w_sum_33_39), .ow_c(w_carry_33_39));
wire w_sum_33_37, w_carry_33_37;
math_adder_carry_save CSA_33_37(.i_a(w_carry_32_50), .i_b(w_carry_32_48), .i_c(w_carry_32_46), .ow_sum(w_sum_33_37), .ow_c(w_carry_33_37));
wire w_sum_33_35, w_carry_33_35;
math_adder_carry_save CSA_33_35(.i_a(w_carry_32_44), .i_b(w_carry_32_42), .i_c(w_carry_32_40), .ow_sum(w_sum_33_35), .ow_c(w_carry_33_35));
wire w_sum_33_33, w_carry_33_33;
math_adder_carry_save CSA_33_33(.i_a(w_carry_32_38), .i_b(w_carry_32_36), .i_c(w_carry_32_34), .ow_sum(w_sum_33_33), .ow_c(w_carry_33_33));
wire w_sum_33_31, w_carry_33_31;
math_adder_carry_save CSA_33_31(.i_a(w_carry_32_32), .i_b(w_carry_32_30), .i_c(w_carry_32_28), .ow_sum(w_sum_33_31), .ow_c(w_carry_33_31));
wire w_sum_33_29, w_carry_33_29;
math_adder_carry_save CSA_33_29(.i_a(w_carry_32_26), .i_b(w_carry_32_24), .i_c(w_carry_32_22), .ow_sum(w_sum_33_29), .ow_c(w_carry_33_29));
wire w_sum_33_27, w_carry_33_27;
math_adder_carry_save CSA_33_27(.i_a(w_carry_32_20), .i_b(w_carry_32_18), .i_c(w_carry_32_16), .ow_sum(w_sum_33_27), .ow_c(w_carry_33_27));
wire w_sum_33_25, w_carry_33_25;
math_adder_carry_save CSA_33_25(.i_a(w_carry_32_14), .i_b(w_carry_32_12), .i_c(w_carry_32_10), .ow_sum(w_sum_33_25), .ow_c(w_carry_33_25));
wire w_sum_33_23, w_carry_33_23;
math_adder_carry_save CSA_33_23(.i_a(w_carry_32_8), .i_b(w_carry_32_6), .i_c(w_carry_32_4), .ow_sum(w_sum_33_23), .ow_c(w_carry_33_23));
wire w_sum_33_21, w_carry_33_21;
math_adder_carry_save CSA_33_21(.i_a(w_carry_32_2), .i_b(w_sum_33_61), .i_c(w_sum_33_59), .ow_sum(w_sum_33_21), .ow_c(w_carry_33_21));
wire w_sum_33_19, w_carry_33_19;
math_adder_carry_save CSA_33_19(.i_a(w_sum_33_57), .i_b(w_sum_33_55), .i_c(w_sum_33_53), .ow_sum(w_sum_33_19), .ow_c(w_carry_33_19));
wire w_sum_33_17, w_carry_33_17;
math_adder_carry_save CSA_33_17(.i_a(w_sum_33_51), .i_b(w_sum_33_49), .i_c(w_sum_33_47), .ow_sum(w_sum_33_17), .ow_c(w_carry_33_17));
wire w_sum_33_15, w_carry_33_15;
math_adder_carry_save CSA_33_15(.i_a(w_sum_33_45), .i_b(w_sum_33_43), .i_c(w_sum_33_41), .ow_sum(w_sum_33_15), .ow_c(w_carry_33_15));
wire w_sum_33_13, w_carry_33_13;
math_adder_carry_save CSA_33_13(.i_a(w_sum_33_39), .i_b(w_sum_33_37), .i_c(w_sum_33_35), .ow_sum(w_sum_33_13), .ow_c(w_carry_33_13));
wire w_sum_33_11, w_carry_33_11;
math_adder_carry_save CSA_33_11(.i_a(w_sum_33_33), .i_b(w_sum_33_31), .i_c(w_sum_33_29), .ow_sum(w_sum_33_11), .ow_c(w_carry_33_11));
wire w_sum_33_9, w_carry_33_9;
math_adder_carry_save CSA_33_9(.i_a(w_sum_33_27), .i_b(w_sum_33_25), .i_c(w_sum_33_23), .ow_sum(w_sum_33_9), .ow_c(w_carry_33_9));
wire w_sum_33_7, w_carry_33_7;
math_adder_carry_save CSA_33_7(.i_a(w_sum_33_21), .i_b(w_sum_33_19), .i_c(w_sum_33_17), .ow_sum(w_sum_33_7), .ow_c(w_carry_33_7));
wire w_sum_33_5, w_carry_33_5;
math_adder_carry_save CSA_33_5(.i_a(w_sum_33_15), .i_b(w_sum_33_13), .i_c(w_sum_33_11), .ow_sum(w_sum_33_5), .ow_c(w_carry_33_5));
wire w_sum_33_3, w_carry_33_3;
math_adder_carry_save CSA_33_3(.i_a(w_sum_33_9), .i_b(w_sum_33_7), .i_c(w_sum_33_5), .ow_sum(w_sum_33_3), .ow_c(w_carry_33_3));
wire w_sum_34_59, w_carry_34_59;
math_adder_carry_save CSA_34_59(.i_a(w_pp_3_31), .i_b(w_pp_4_30), .i_c(w_pp_5_29), .ow_sum(w_sum_34_59), .ow_c(w_carry_34_59));
wire w_sum_34_57, w_carry_34_57;
math_adder_carry_save CSA_34_57(.i_a(w_pp_6_28), .i_b(w_pp_7_27), .i_c(w_pp_8_26), .ow_sum(w_sum_34_57), .ow_c(w_carry_34_57));
wire w_sum_34_55, w_carry_34_55;
math_adder_carry_save CSA_34_55(.i_a(w_pp_9_25), .i_b(w_pp_10_24), .i_c(w_pp_11_23), .ow_sum(w_sum_34_55), .ow_c(w_carry_34_55));
wire w_sum_34_53, w_carry_34_53;
math_adder_carry_save CSA_34_53(.i_a(w_pp_12_22), .i_b(w_pp_13_21), .i_c(w_pp_14_20), .ow_sum(w_sum_34_53), .ow_c(w_carry_34_53));
wire w_sum_34_51, w_carry_34_51;
math_adder_carry_save CSA_34_51(.i_a(w_pp_15_19), .i_b(w_pp_16_18), .i_c(w_pp_17_17), .ow_sum(w_sum_34_51), .ow_c(w_carry_34_51));
wire w_sum_34_49, w_carry_34_49;
math_adder_carry_save CSA_34_49(.i_a(w_pp_18_16), .i_b(w_pp_19_15), .i_c(w_pp_20_14), .ow_sum(w_sum_34_49), .ow_c(w_carry_34_49));
wire w_sum_34_47, w_carry_34_47;
math_adder_carry_save CSA_34_47(.i_a(w_pp_21_13), .i_b(w_pp_22_12), .i_c(w_pp_23_11), .ow_sum(w_sum_34_47), .ow_c(w_carry_34_47));
wire w_sum_34_45, w_carry_34_45;
math_adder_carry_save CSA_34_45(.i_a(w_pp_24_10), .i_b(w_pp_25_9), .i_c(w_pp_26_8), .ow_sum(w_sum_34_45), .ow_c(w_carry_34_45));
wire w_sum_34_43, w_carry_34_43;
math_adder_carry_save CSA_34_43(.i_a(w_pp_27_7), .i_b(w_pp_28_6), .i_c(w_pp_29_5), .ow_sum(w_sum_34_43), .ow_c(w_carry_34_43));
wire w_sum_34_41, w_carry_34_41;
math_adder_carry_save CSA_34_41(.i_a(w_pp_30_4), .i_b(w_pp_31_3), .i_c(w_carry_33_61), .ow_sum(w_sum_34_41), .ow_c(w_carry_34_41));
wire w_sum_34_39, w_carry_34_39;
math_adder_carry_save CSA_34_39(.i_a(w_carry_33_59), .i_b(w_carry_33_57), .i_c(w_carry_33_55), .ow_sum(w_sum_34_39), .ow_c(w_carry_34_39));
wire w_sum_34_37, w_carry_34_37;
math_adder_carry_save CSA_34_37(.i_a(w_carry_33_53), .i_b(w_carry_33_51), .i_c(w_carry_33_49), .ow_sum(w_sum_34_37), .ow_c(w_carry_34_37));
wire w_sum_34_35, w_carry_34_35;
math_adder_carry_save CSA_34_35(.i_a(w_carry_33_47), .i_b(w_carry_33_45), .i_c(w_carry_33_43), .ow_sum(w_sum_34_35), .ow_c(w_carry_34_35));
wire w_sum_34_33, w_carry_34_33;
math_adder_carry_save CSA_34_33(.i_a(w_carry_33_41), .i_b(w_carry_33_39), .i_c(w_carry_33_37), .ow_sum(w_sum_34_33), .ow_c(w_carry_34_33));
wire w_sum_34_31, w_carry_34_31;
math_adder_carry_save CSA_34_31(.i_a(w_carry_33_35), .i_b(w_carry_33_33), .i_c(w_carry_33_31), .ow_sum(w_sum_34_31), .ow_c(w_carry_34_31));
wire w_sum_34_29, w_carry_34_29;
math_adder_carry_save CSA_34_29(.i_a(w_carry_33_29), .i_b(w_carry_33_27), .i_c(w_carry_33_25), .ow_sum(w_sum_34_29), .ow_c(w_carry_34_29));
wire w_sum_34_27, w_carry_34_27;
math_adder_carry_save CSA_34_27(.i_a(w_carry_33_23), .i_b(w_carry_33_21), .i_c(w_carry_33_19), .ow_sum(w_sum_34_27), .ow_c(w_carry_34_27));
wire w_sum_34_25, w_carry_34_25;
math_adder_carry_save CSA_34_25(.i_a(w_carry_33_17), .i_b(w_carry_33_15), .i_c(w_carry_33_13), .ow_sum(w_sum_34_25), .ow_c(w_carry_34_25));
wire w_sum_34_23, w_carry_34_23;
math_adder_carry_save CSA_34_23(.i_a(w_carry_33_11), .i_b(w_carry_33_9), .i_c(w_carry_33_7), .ow_sum(w_sum_34_23), .ow_c(w_carry_34_23));
wire w_sum_34_21, w_carry_34_21;
math_adder_carry_save CSA_34_21(.i_a(w_carry_33_5), .i_b(w_carry_33_3), .i_c(w_sum_34_59), .ow_sum(w_sum_34_21), .ow_c(w_carry_34_21));
wire w_sum_34_19, w_carry_34_19;
math_adder_carry_save CSA_34_19(.i_a(w_sum_34_57), .i_b(w_sum_34_55), .i_c(w_sum_34_53), .ow_sum(w_sum_34_19), .ow_c(w_carry_34_19));
wire w_sum_34_17, w_carry_34_17;
math_adder_carry_save CSA_34_17(.i_a(w_sum_34_51), .i_b(w_sum_34_49), .i_c(w_sum_34_47), .ow_sum(w_sum_34_17), .ow_c(w_carry_34_17));
wire w_sum_34_15, w_carry_34_15;
math_adder_carry_save CSA_34_15(.i_a(w_sum_34_45), .i_b(w_sum_34_43), .i_c(w_sum_34_41), .ow_sum(w_sum_34_15), .ow_c(w_carry_34_15));
wire w_sum_34_13, w_carry_34_13;
math_adder_carry_save CSA_34_13(.i_a(w_sum_34_39), .i_b(w_sum_34_37), .i_c(w_sum_34_35), .ow_sum(w_sum_34_13), .ow_c(w_carry_34_13));
wire w_sum_34_11, w_carry_34_11;
math_adder_carry_save CSA_34_11(.i_a(w_sum_34_33), .i_b(w_sum_34_31), .i_c(w_sum_34_29), .ow_sum(w_sum_34_11), .ow_c(w_carry_34_11));
wire w_sum_34_9, w_carry_34_9;
math_adder_carry_save CSA_34_9(.i_a(w_sum_34_27), .i_b(w_sum_34_25), .i_c(w_sum_34_23), .ow_sum(w_sum_34_9), .ow_c(w_carry_34_9));
wire w_sum_34_7, w_carry_34_7;
math_adder_carry_save CSA_34_7(.i_a(w_sum_34_21), .i_b(w_sum_34_19), .i_c(w_sum_34_17), .ow_sum(w_sum_34_7), .ow_c(w_carry_34_7));
wire w_sum_34_5, w_carry_34_5;
math_adder_carry_save CSA_34_5(.i_a(w_sum_34_15), .i_b(w_sum_34_13), .i_c(w_sum_34_11), .ow_sum(w_sum_34_5), .ow_c(w_carry_34_5));
wire w_sum_34_3, w_carry_34_3;
math_adder_carry_save CSA_34_3(.i_a(w_sum_34_9), .i_b(w_sum_34_7), .i_c(w_sum_34_5), .ow_sum(w_sum_34_3), .ow_c(w_carry_34_3));
wire w_sum_35_57, w_carry_35_57;
math_adder_carry_save CSA_35_57(.i_a(w_pp_4_31), .i_b(w_pp_5_30), .i_c(w_pp_6_29), .ow_sum(w_sum_35_57), .ow_c(w_carry_35_57));
wire w_sum_35_55, w_carry_35_55;
math_adder_carry_save CSA_35_55(.i_a(w_pp_7_28), .i_b(w_pp_8_27), .i_c(w_pp_9_26), .ow_sum(w_sum_35_55), .ow_c(w_carry_35_55));
wire w_sum_35_53, w_carry_35_53;
math_adder_carry_save CSA_35_53(.i_a(w_pp_10_25), .i_b(w_pp_11_24), .i_c(w_pp_12_23), .ow_sum(w_sum_35_53), .ow_c(w_carry_35_53));
wire w_sum_35_51, w_carry_35_51;
math_adder_carry_save CSA_35_51(.i_a(w_pp_13_22), .i_b(w_pp_14_21), .i_c(w_pp_15_20), .ow_sum(w_sum_35_51), .ow_c(w_carry_35_51));
wire w_sum_35_49, w_carry_35_49;
math_adder_carry_save CSA_35_49(.i_a(w_pp_16_19), .i_b(w_pp_17_18), .i_c(w_pp_18_17), .ow_sum(w_sum_35_49), .ow_c(w_carry_35_49));
wire w_sum_35_47, w_carry_35_47;
math_adder_carry_save CSA_35_47(.i_a(w_pp_19_16), .i_b(w_pp_20_15), .i_c(w_pp_21_14), .ow_sum(w_sum_35_47), .ow_c(w_carry_35_47));
wire w_sum_35_45, w_carry_35_45;
math_adder_carry_save CSA_35_45(.i_a(w_pp_22_13), .i_b(w_pp_23_12), .i_c(w_pp_24_11), .ow_sum(w_sum_35_45), .ow_c(w_carry_35_45));
wire w_sum_35_43, w_carry_35_43;
math_adder_carry_save CSA_35_43(.i_a(w_pp_25_10), .i_b(w_pp_26_9), .i_c(w_pp_27_8), .ow_sum(w_sum_35_43), .ow_c(w_carry_35_43));
wire w_sum_35_41, w_carry_35_41;
math_adder_carry_save CSA_35_41(.i_a(w_pp_28_7), .i_b(w_pp_29_6), .i_c(w_pp_30_5), .ow_sum(w_sum_35_41), .ow_c(w_carry_35_41));
wire w_sum_35_39, w_carry_35_39;
math_adder_carry_save CSA_35_39(.i_a(w_pp_31_4), .i_b(w_carry_34_59), .i_c(w_carry_34_57), .ow_sum(w_sum_35_39), .ow_c(w_carry_35_39));
wire w_sum_35_37, w_carry_35_37;
math_adder_carry_save CSA_35_37(.i_a(w_carry_34_55), .i_b(w_carry_34_53), .i_c(w_carry_34_51), .ow_sum(w_sum_35_37), .ow_c(w_carry_35_37));
wire w_sum_35_35, w_carry_35_35;
math_adder_carry_save CSA_35_35(.i_a(w_carry_34_49), .i_b(w_carry_34_47), .i_c(w_carry_34_45), .ow_sum(w_sum_35_35), .ow_c(w_carry_35_35));
wire w_sum_35_33, w_carry_35_33;
math_adder_carry_save CSA_35_33(.i_a(w_carry_34_43), .i_b(w_carry_34_41), .i_c(w_carry_34_39), .ow_sum(w_sum_35_33), .ow_c(w_carry_35_33));
wire w_sum_35_31, w_carry_35_31;
math_adder_carry_save CSA_35_31(.i_a(w_carry_34_37), .i_b(w_carry_34_35), .i_c(w_carry_34_33), .ow_sum(w_sum_35_31), .ow_c(w_carry_35_31));
wire w_sum_35_29, w_carry_35_29;
math_adder_carry_save CSA_35_29(.i_a(w_carry_34_31), .i_b(w_carry_34_29), .i_c(w_carry_34_27), .ow_sum(w_sum_35_29), .ow_c(w_carry_35_29));
wire w_sum_35_27, w_carry_35_27;
math_adder_carry_save CSA_35_27(.i_a(w_carry_34_25), .i_b(w_carry_34_23), .i_c(w_carry_34_21), .ow_sum(w_sum_35_27), .ow_c(w_carry_35_27));
wire w_sum_35_25, w_carry_35_25;
math_adder_carry_save CSA_35_25(.i_a(w_carry_34_19), .i_b(w_carry_34_17), .i_c(w_carry_34_15), .ow_sum(w_sum_35_25), .ow_c(w_carry_35_25));
wire w_sum_35_23, w_carry_35_23;
math_adder_carry_save CSA_35_23(.i_a(w_carry_34_13), .i_b(w_carry_34_11), .i_c(w_carry_34_9), .ow_sum(w_sum_35_23), .ow_c(w_carry_35_23));
wire w_sum_35_21, w_carry_35_21;
math_adder_carry_save CSA_35_21(.i_a(w_carry_34_7), .i_b(w_carry_34_5), .i_c(w_carry_34_3), .ow_sum(w_sum_35_21), .ow_c(w_carry_35_21));
wire w_sum_35_19, w_carry_35_19;
math_adder_carry_save CSA_35_19(.i_a(w_sum_35_57), .i_b(w_sum_35_55), .i_c(w_sum_35_53), .ow_sum(w_sum_35_19), .ow_c(w_carry_35_19));
wire w_sum_35_17, w_carry_35_17;
math_adder_carry_save CSA_35_17(.i_a(w_sum_35_51), .i_b(w_sum_35_49), .i_c(w_sum_35_47), .ow_sum(w_sum_35_17), .ow_c(w_carry_35_17));
wire w_sum_35_15, w_carry_35_15;
math_adder_carry_save CSA_35_15(.i_a(w_sum_35_45), .i_b(w_sum_35_43), .i_c(w_sum_35_41), .ow_sum(w_sum_35_15), .ow_c(w_carry_35_15));
wire w_sum_35_13, w_carry_35_13;
math_adder_carry_save CSA_35_13(.i_a(w_sum_35_39), .i_b(w_sum_35_37), .i_c(w_sum_35_35), .ow_sum(w_sum_35_13), .ow_c(w_carry_35_13));
wire w_sum_35_11, w_carry_35_11;
math_adder_carry_save CSA_35_11(.i_a(w_sum_35_33), .i_b(w_sum_35_31), .i_c(w_sum_35_29), .ow_sum(w_sum_35_11), .ow_c(w_carry_35_11));
wire w_sum_35_9, w_carry_35_9;
math_adder_carry_save CSA_35_9(.i_a(w_sum_35_27), .i_b(w_sum_35_25), .i_c(w_sum_35_23), .ow_sum(w_sum_35_9), .ow_c(w_carry_35_9));
wire w_sum_35_7, w_carry_35_7;
math_adder_carry_save CSA_35_7(.i_a(w_sum_35_21), .i_b(w_sum_35_19), .i_c(w_sum_35_17), .ow_sum(w_sum_35_7), .ow_c(w_carry_35_7));
wire w_sum_35_5, w_carry_35_5;
math_adder_carry_save CSA_35_5(.i_a(w_sum_35_15), .i_b(w_sum_35_13), .i_c(w_sum_35_11), .ow_sum(w_sum_35_5), .ow_c(w_carry_35_5));
wire w_sum_35_3, w_carry_35_3;
math_adder_carry_save CSA_35_3(.i_a(w_sum_35_9), .i_b(w_sum_35_7), .i_c(w_sum_35_5), .ow_sum(w_sum_35_3), .ow_c(w_carry_35_3));
wire w_sum_36_55, w_carry_36_55;
math_adder_carry_save CSA_36_55(.i_a(w_pp_5_31), .i_b(w_pp_6_30), .i_c(w_pp_7_29), .ow_sum(w_sum_36_55), .ow_c(w_carry_36_55));
wire w_sum_36_53, w_carry_36_53;
math_adder_carry_save CSA_36_53(.i_a(w_pp_8_28), .i_b(w_pp_9_27), .i_c(w_pp_10_26), .ow_sum(w_sum_36_53), .ow_c(w_carry_36_53));
wire w_sum_36_51, w_carry_36_51;
math_adder_carry_save CSA_36_51(.i_a(w_pp_11_25), .i_b(w_pp_12_24), .i_c(w_pp_13_23), .ow_sum(w_sum_36_51), .ow_c(w_carry_36_51));
wire w_sum_36_49, w_carry_36_49;
math_adder_carry_save CSA_36_49(.i_a(w_pp_14_22), .i_b(w_pp_15_21), .i_c(w_pp_16_20), .ow_sum(w_sum_36_49), .ow_c(w_carry_36_49));
wire w_sum_36_47, w_carry_36_47;
math_adder_carry_save CSA_36_47(.i_a(w_pp_17_19), .i_b(w_pp_18_18), .i_c(w_pp_19_17), .ow_sum(w_sum_36_47), .ow_c(w_carry_36_47));
wire w_sum_36_45, w_carry_36_45;
math_adder_carry_save CSA_36_45(.i_a(w_pp_20_16), .i_b(w_pp_21_15), .i_c(w_pp_22_14), .ow_sum(w_sum_36_45), .ow_c(w_carry_36_45));
wire w_sum_36_43, w_carry_36_43;
math_adder_carry_save CSA_36_43(.i_a(w_pp_23_13), .i_b(w_pp_24_12), .i_c(w_pp_25_11), .ow_sum(w_sum_36_43), .ow_c(w_carry_36_43));
wire w_sum_36_41, w_carry_36_41;
math_adder_carry_save CSA_36_41(.i_a(w_pp_26_10), .i_b(w_pp_27_9), .i_c(w_pp_28_8), .ow_sum(w_sum_36_41), .ow_c(w_carry_36_41));
wire w_sum_36_39, w_carry_36_39;
math_adder_carry_save CSA_36_39(.i_a(w_pp_29_7), .i_b(w_pp_30_6), .i_c(w_pp_31_5), .ow_sum(w_sum_36_39), .ow_c(w_carry_36_39));
wire w_sum_36_37, w_carry_36_37;
math_adder_carry_save CSA_36_37(.i_a(w_carry_35_57), .i_b(w_carry_35_55), .i_c(w_carry_35_53), .ow_sum(w_sum_36_37), .ow_c(w_carry_36_37));
wire w_sum_36_35, w_carry_36_35;
math_adder_carry_save CSA_36_35(.i_a(w_carry_35_51), .i_b(w_carry_35_49), .i_c(w_carry_35_47), .ow_sum(w_sum_36_35), .ow_c(w_carry_36_35));
wire w_sum_36_33, w_carry_36_33;
math_adder_carry_save CSA_36_33(.i_a(w_carry_35_45), .i_b(w_carry_35_43), .i_c(w_carry_35_41), .ow_sum(w_sum_36_33), .ow_c(w_carry_36_33));
wire w_sum_36_31, w_carry_36_31;
math_adder_carry_save CSA_36_31(.i_a(w_carry_35_39), .i_b(w_carry_35_37), .i_c(w_carry_35_35), .ow_sum(w_sum_36_31), .ow_c(w_carry_36_31));
wire w_sum_36_29, w_carry_36_29;
math_adder_carry_save CSA_36_29(.i_a(w_carry_35_33), .i_b(w_carry_35_31), .i_c(w_carry_35_29), .ow_sum(w_sum_36_29), .ow_c(w_carry_36_29));
wire w_sum_36_27, w_carry_36_27;
math_adder_carry_save CSA_36_27(.i_a(w_carry_35_27), .i_b(w_carry_35_25), .i_c(w_carry_35_23), .ow_sum(w_sum_36_27), .ow_c(w_carry_36_27));
wire w_sum_36_25, w_carry_36_25;
math_adder_carry_save CSA_36_25(.i_a(w_carry_35_21), .i_b(w_carry_35_19), .i_c(w_carry_35_17), .ow_sum(w_sum_36_25), .ow_c(w_carry_36_25));
wire w_sum_36_23, w_carry_36_23;
math_adder_carry_save CSA_36_23(.i_a(w_carry_35_15), .i_b(w_carry_35_13), .i_c(w_carry_35_11), .ow_sum(w_sum_36_23), .ow_c(w_carry_36_23));
wire w_sum_36_21, w_carry_36_21;
math_adder_carry_save CSA_36_21(.i_a(w_carry_35_9), .i_b(w_carry_35_7), .i_c(w_carry_35_5), .ow_sum(w_sum_36_21), .ow_c(w_carry_36_21));
wire w_sum_36_19, w_carry_36_19;
math_adder_carry_save CSA_36_19(.i_a(w_carry_35_3), .i_b(w_sum_36_55), .i_c(w_sum_36_53), .ow_sum(w_sum_36_19), .ow_c(w_carry_36_19));
wire w_sum_36_17, w_carry_36_17;
math_adder_carry_save CSA_36_17(.i_a(w_sum_36_51), .i_b(w_sum_36_49), .i_c(w_sum_36_47), .ow_sum(w_sum_36_17), .ow_c(w_carry_36_17));
wire w_sum_36_15, w_carry_36_15;
math_adder_carry_save CSA_36_15(.i_a(w_sum_36_45), .i_b(w_sum_36_43), .i_c(w_sum_36_41), .ow_sum(w_sum_36_15), .ow_c(w_carry_36_15));
wire w_sum_36_13, w_carry_36_13;
math_adder_carry_save CSA_36_13(.i_a(w_sum_36_39), .i_b(w_sum_36_37), .i_c(w_sum_36_35), .ow_sum(w_sum_36_13), .ow_c(w_carry_36_13));
wire w_sum_36_11, w_carry_36_11;
math_adder_carry_save CSA_36_11(.i_a(w_sum_36_33), .i_b(w_sum_36_31), .i_c(w_sum_36_29), .ow_sum(w_sum_36_11), .ow_c(w_carry_36_11));
wire w_sum_36_9, w_carry_36_9;
math_adder_carry_save CSA_36_9(.i_a(w_sum_36_27), .i_b(w_sum_36_25), .i_c(w_sum_36_23), .ow_sum(w_sum_36_9), .ow_c(w_carry_36_9));
wire w_sum_36_7, w_carry_36_7;
math_adder_carry_save CSA_36_7(.i_a(w_sum_36_21), .i_b(w_sum_36_19), .i_c(w_sum_36_17), .ow_sum(w_sum_36_7), .ow_c(w_carry_36_7));
wire w_sum_36_5, w_carry_36_5;
math_adder_carry_save CSA_36_5(.i_a(w_sum_36_15), .i_b(w_sum_36_13), .i_c(w_sum_36_11), .ow_sum(w_sum_36_5), .ow_c(w_carry_36_5));
wire w_sum_36_3, w_carry_36_3;
math_adder_carry_save CSA_36_3(.i_a(w_sum_36_9), .i_b(w_sum_36_7), .i_c(w_sum_36_5), .ow_sum(w_sum_36_3), .ow_c(w_carry_36_3));
wire w_sum_37_53, w_carry_37_53;
math_adder_carry_save CSA_37_53(.i_a(w_pp_6_31), .i_b(w_pp_7_30), .i_c(w_pp_8_29), .ow_sum(w_sum_37_53), .ow_c(w_carry_37_53));
wire w_sum_37_51, w_carry_37_51;
math_adder_carry_save CSA_37_51(.i_a(w_pp_9_28), .i_b(w_pp_10_27), .i_c(w_pp_11_26), .ow_sum(w_sum_37_51), .ow_c(w_carry_37_51));
wire w_sum_37_49, w_carry_37_49;
math_adder_carry_save CSA_37_49(.i_a(w_pp_12_25), .i_b(w_pp_13_24), .i_c(w_pp_14_23), .ow_sum(w_sum_37_49), .ow_c(w_carry_37_49));
wire w_sum_37_47, w_carry_37_47;
math_adder_carry_save CSA_37_47(.i_a(w_pp_15_22), .i_b(w_pp_16_21), .i_c(w_pp_17_20), .ow_sum(w_sum_37_47), .ow_c(w_carry_37_47));
wire w_sum_37_45, w_carry_37_45;
math_adder_carry_save CSA_37_45(.i_a(w_pp_18_19), .i_b(w_pp_19_18), .i_c(w_pp_20_17), .ow_sum(w_sum_37_45), .ow_c(w_carry_37_45));
wire w_sum_37_43, w_carry_37_43;
math_adder_carry_save CSA_37_43(.i_a(w_pp_21_16), .i_b(w_pp_22_15), .i_c(w_pp_23_14), .ow_sum(w_sum_37_43), .ow_c(w_carry_37_43));
wire w_sum_37_41, w_carry_37_41;
math_adder_carry_save CSA_37_41(.i_a(w_pp_24_13), .i_b(w_pp_25_12), .i_c(w_pp_26_11), .ow_sum(w_sum_37_41), .ow_c(w_carry_37_41));
wire w_sum_37_39, w_carry_37_39;
math_adder_carry_save CSA_37_39(.i_a(w_pp_27_10), .i_b(w_pp_28_9), .i_c(w_pp_29_8), .ow_sum(w_sum_37_39), .ow_c(w_carry_37_39));
wire w_sum_37_37, w_carry_37_37;
math_adder_carry_save CSA_37_37(.i_a(w_pp_30_7), .i_b(w_pp_31_6), .i_c(w_carry_36_55), .ow_sum(w_sum_37_37), .ow_c(w_carry_37_37));
wire w_sum_37_35, w_carry_37_35;
math_adder_carry_save CSA_37_35(.i_a(w_carry_36_53), .i_b(w_carry_36_51), .i_c(w_carry_36_49), .ow_sum(w_sum_37_35), .ow_c(w_carry_37_35));
wire w_sum_37_33, w_carry_37_33;
math_adder_carry_save CSA_37_33(.i_a(w_carry_36_47), .i_b(w_carry_36_45), .i_c(w_carry_36_43), .ow_sum(w_sum_37_33), .ow_c(w_carry_37_33));
wire w_sum_37_31, w_carry_37_31;
math_adder_carry_save CSA_37_31(.i_a(w_carry_36_41), .i_b(w_carry_36_39), .i_c(w_carry_36_37), .ow_sum(w_sum_37_31), .ow_c(w_carry_37_31));
wire w_sum_37_29, w_carry_37_29;
math_adder_carry_save CSA_37_29(.i_a(w_carry_36_35), .i_b(w_carry_36_33), .i_c(w_carry_36_31), .ow_sum(w_sum_37_29), .ow_c(w_carry_37_29));
wire w_sum_37_27, w_carry_37_27;
math_adder_carry_save CSA_37_27(.i_a(w_carry_36_29), .i_b(w_carry_36_27), .i_c(w_carry_36_25), .ow_sum(w_sum_37_27), .ow_c(w_carry_37_27));
wire w_sum_37_25, w_carry_37_25;
math_adder_carry_save CSA_37_25(.i_a(w_carry_36_23), .i_b(w_carry_36_21), .i_c(w_carry_36_19), .ow_sum(w_sum_37_25), .ow_c(w_carry_37_25));
wire w_sum_37_23, w_carry_37_23;
math_adder_carry_save CSA_37_23(.i_a(w_carry_36_17), .i_b(w_carry_36_15), .i_c(w_carry_36_13), .ow_sum(w_sum_37_23), .ow_c(w_carry_37_23));
wire w_sum_37_21, w_carry_37_21;
math_adder_carry_save CSA_37_21(.i_a(w_carry_36_11), .i_b(w_carry_36_9), .i_c(w_carry_36_7), .ow_sum(w_sum_37_21), .ow_c(w_carry_37_21));
wire w_sum_37_19, w_carry_37_19;
math_adder_carry_save CSA_37_19(.i_a(w_carry_36_5), .i_b(w_carry_36_3), .i_c(w_sum_37_53), .ow_sum(w_sum_37_19), .ow_c(w_carry_37_19));
wire w_sum_37_17, w_carry_37_17;
math_adder_carry_save CSA_37_17(.i_a(w_sum_37_51), .i_b(w_sum_37_49), .i_c(w_sum_37_47), .ow_sum(w_sum_37_17), .ow_c(w_carry_37_17));
wire w_sum_37_15, w_carry_37_15;
math_adder_carry_save CSA_37_15(.i_a(w_sum_37_45), .i_b(w_sum_37_43), .i_c(w_sum_37_41), .ow_sum(w_sum_37_15), .ow_c(w_carry_37_15));
wire w_sum_37_13, w_carry_37_13;
math_adder_carry_save CSA_37_13(.i_a(w_sum_37_39), .i_b(w_sum_37_37), .i_c(w_sum_37_35), .ow_sum(w_sum_37_13), .ow_c(w_carry_37_13));
wire w_sum_37_11, w_carry_37_11;
math_adder_carry_save CSA_37_11(.i_a(w_sum_37_33), .i_b(w_sum_37_31), .i_c(w_sum_37_29), .ow_sum(w_sum_37_11), .ow_c(w_carry_37_11));
wire w_sum_37_9, w_carry_37_9;
math_adder_carry_save CSA_37_9(.i_a(w_sum_37_27), .i_b(w_sum_37_25), .i_c(w_sum_37_23), .ow_sum(w_sum_37_9), .ow_c(w_carry_37_9));
wire w_sum_37_7, w_carry_37_7;
math_adder_carry_save CSA_37_7(.i_a(w_sum_37_21), .i_b(w_sum_37_19), .i_c(w_sum_37_17), .ow_sum(w_sum_37_7), .ow_c(w_carry_37_7));
wire w_sum_37_5, w_carry_37_5;
math_adder_carry_save CSA_37_5(.i_a(w_sum_37_15), .i_b(w_sum_37_13), .i_c(w_sum_37_11), .ow_sum(w_sum_37_5), .ow_c(w_carry_37_5));
wire w_sum_37_3, w_carry_37_3;
math_adder_carry_save CSA_37_3(.i_a(w_sum_37_9), .i_b(w_sum_37_7), .i_c(w_sum_37_5), .ow_sum(w_sum_37_3), .ow_c(w_carry_37_3));
wire w_sum_38_51, w_carry_38_51;
math_adder_carry_save CSA_38_51(.i_a(w_pp_7_31), .i_b(w_pp_8_30), .i_c(w_pp_9_29), .ow_sum(w_sum_38_51), .ow_c(w_carry_38_51));
wire w_sum_38_49, w_carry_38_49;
math_adder_carry_save CSA_38_49(.i_a(w_pp_10_28), .i_b(w_pp_11_27), .i_c(w_pp_12_26), .ow_sum(w_sum_38_49), .ow_c(w_carry_38_49));
wire w_sum_38_47, w_carry_38_47;
math_adder_carry_save CSA_38_47(.i_a(w_pp_13_25), .i_b(w_pp_14_24), .i_c(w_pp_15_23), .ow_sum(w_sum_38_47), .ow_c(w_carry_38_47));
wire w_sum_38_45, w_carry_38_45;
math_adder_carry_save CSA_38_45(.i_a(w_pp_16_22), .i_b(w_pp_17_21), .i_c(w_pp_18_20), .ow_sum(w_sum_38_45), .ow_c(w_carry_38_45));
wire w_sum_38_43, w_carry_38_43;
math_adder_carry_save CSA_38_43(.i_a(w_pp_19_19), .i_b(w_pp_20_18), .i_c(w_pp_21_17), .ow_sum(w_sum_38_43), .ow_c(w_carry_38_43));
wire w_sum_38_41, w_carry_38_41;
math_adder_carry_save CSA_38_41(.i_a(w_pp_22_16), .i_b(w_pp_23_15), .i_c(w_pp_24_14), .ow_sum(w_sum_38_41), .ow_c(w_carry_38_41));
wire w_sum_38_39, w_carry_38_39;
math_adder_carry_save CSA_38_39(.i_a(w_pp_25_13), .i_b(w_pp_26_12), .i_c(w_pp_27_11), .ow_sum(w_sum_38_39), .ow_c(w_carry_38_39));
wire w_sum_38_37, w_carry_38_37;
math_adder_carry_save CSA_38_37(.i_a(w_pp_28_10), .i_b(w_pp_29_9), .i_c(w_pp_30_8), .ow_sum(w_sum_38_37), .ow_c(w_carry_38_37));
wire w_sum_38_35, w_carry_38_35;
math_adder_carry_save CSA_38_35(.i_a(w_pp_31_7), .i_b(w_carry_37_53), .i_c(w_carry_37_51), .ow_sum(w_sum_38_35), .ow_c(w_carry_38_35));
wire w_sum_38_33, w_carry_38_33;
math_adder_carry_save CSA_38_33(.i_a(w_carry_37_49), .i_b(w_carry_37_47), .i_c(w_carry_37_45), .ow_sum(w_sum_38_33), .ow_c(w_carry_38_33));
wire w_sum_38_31, w_carry_38_31;
math_adder_carry_save CSA_38_31(.i_a(w_carry_37_43), .i_b(w_carry_37_41), .i_c(w_carry_37_39), .ow_sum(w_sum_38_31), .ow_c(w_carry_38_31));
wire w_sum_38_29, w_carry_38_29;
math_adder_carry_save CSA_38_29(.i_a(w_carry_37_37), .i_b(w_carry_37_35), .i_c(w_carry_37_33), .ow_sum(w_sum_38_29), .ow_c(w_carry_38_29));
wire w_sum_38_27, w_carry_38_27;
math_adder_carry_save CSA_38_27(.i_a(w_carry_37_31), .i_b(w_carry_37_29), .i_c(w_carry_37_27), .ow_sum(w_sum_38_27), .ow_c(w_carry_38_27));
wire w_sum_38_25, w_carry_38_25;
math_adder_carry_save CSA_38_25(.i_a(w_carry_37_25), .i_b(w_carry_37_23), .i_c(w_carry_37_21), .ow_sum(w_sum_38_25), .ow_c(w_carry_38_25));
wire w_sum_38_23, w_carry_38_23;
math_adder_carry_save CSA_38_23(.i_a(w_carry_37_19), .i_b(w_carry_37_17), .i_c(w_carry_37_15), .ow_sum(w_sum_38_23), .ow_c(w_carry_38_23));
wire w_sum_38_21, w_carry_38_21;
math_adder_carry_save CSA_38_21(.i_a(w_carry_37_13), .i_b(w_carry_37_11), .i_c(w_carry_37_9), .ow_sum(w_sum_38_21), .ow_c(w_carry_38_21));
wire w_sum_38_19, w_carry_38_19;
math_adder_carry_save CSA_38_19(.i_a(w_carry_37_7), .i_b(w_carry_37_5), .i_c(w_carry_37_3), .ow_sum(w_sum_38_19), .ow_c(w_carry_38_19));
wire w_sum_38_17, w_carry_38_17;
math_adder_carry_save CSA_38_17(.i_a(w_sum_38_51), .i_b(w_sum_38_49), .i_c(w_sum_38_47), .ow_sum(w_sum_38_17), .ow_c(w_carry_38_17));
wire w_sum_38_15, w_carry_38_15;
math_adder_carry_save CSA_38_15(.i_a(w_sum_38_45), .i_b(w_sum_38_43), .i_c(w_sum_38_41), .ow_sum(w_sum_38_15), .ow_c(w_carry_38_15));
wire w_sum_38_13, w_carry_38_13;
math_adder_carry_save CSA_38_13(.i_a(w_sum_38_39), .i_b(w_sum_38_37), .i_c(w_sum_38_35), .ow_sum(w_sum_38_13), .ow_c(w_carry_38_13));
wire w_sum_38_11, w_carry_38_11;
math_adder_carry_save CSA_38_11(.i_a(w_sum_38_33), .i_b(w_sum_38_31), .i_c(w_sum_38_29), .ow_sum(w_sum_38_11), .ow_c(w_carry_38_11));
wire w_sum_38_9, w_carry_38_9;
math_adder_carry_save CSA_38_9(.i_a(w_sum_38_27), .i_b(w_sum_38_25), .i_c(w_sum_38_23), .ow_sum(w_sum_38_9), .ow_c(w_carry_38_9));
wire w_sum_38_7, w_carry_38_7;
math_adder_carry_save CSA_38_7(.i_a(w_sum_38_21), .i_b(w_sum_38_19), .i_c(w_sum_38_17), .ow_sum(w_sum_38_7), .ow_c(w_carry_38_7));
wire w_sum_38_5, w_carry_38_5;
math_adder_carry_save CSA_38_5(.i_a(w_sum_38_15), .i_b(w_sum_38_13), .i_c(w_sum_38_11), .ow_sum(w_sum_38_5), .ow_c(w_carry_38_5));
wire w_sum_38_3, w_carry_38_3;
math_adder_carry_save CSA_38_3(.i_a(w_sum_38_9), .i_b(w_sum_38_7), .i_c(w_sum_38_5), .ow_sum(w_sum_38_3), .ow_c(w_carry_38_3));
wire w_sum_39_49, w_carry_39_49;
math_adder_carry_save CSA_39_49(.i_a(w_pp_8_31), .i_b(w_pp_9_30), .i_c(w_pp_10_29), .ow_sum(w_sum_39_49), .ow_c(w_carry_39_49));
wire w_sum_39_47, w_carry_39_47;
math_adder_carry_save CSA_39_47(.i_a(w_pp_11_28), .i_b(w_pp_12_27), .i_c(w_pp_13_26), .ow_sum(w_sum_39_47), .ow_c(w_carry_39_47));
wire w_sum_39_45, w_carry_39_45;
math_adder_carry_save CSA_39_45(.i_a(w_pp_14_25), .i_b(w_pp_15_24), .i_c(w_pp_16_23), .ow_sum(w_sum_39_45), .ow_c(w_carry_39_45));
wire w_sum_39_43, w_carry_39_43;
math_adder_carry_save CSA_39_43(.i_a(w_pp_17_22), .i_b(w_pp_18_21), .i_c(w_pp_19_20), .ow_sum(w_sum_39_43), .ow_c(w_carry_39_43));
wire w_sum_39_41, w_carry_39_41;
math_adder_carry_save CSA_39_41(.i_a(w_pp_20_19), .i_b(w_pp_21_18), .i_c(w_pp_22_17), .ow_sum(w_sum_39_41), .ow_c(w_carry_39_41));
wire w_sum_39_39, w_carry_39_39;
math_adder_carry_save CSA_39_39(.i_a(w_pp_23_16), .i_b(w_pp_24_15), .i_c(w_pp_25_14), .ow_sum(w_sum_39_39), .ow_c(w_carry_39_39));
wire w_sum_39_37, w_carry_39_37;
math_adder_carry_save CSA_39_37(.i_a(w_pp_26_13), .i_b(w_pp_27_12), .i_c(w_pp_28_11), .ow_sum(w_sum_39_37), .ow_c(w_carry_39_37));
wire w_sum_39_35, w_carry_39_35;
math_adder_carry_save CSA_39_35(.i_a(w_pp_29_10), .i_b(w_pp_30_9), .i_c(w_pp_31_8), .ow_sum(w_sum_39_35), .ow_c(w_carry_39_35));
wire w_sum_39_33, w_carry_39_33;
math_adder_carry_save CSA_39_33(.i_a(w_carry_38_51), .i_b(w_carry_38_49), .i_c(w_carry_38_47), .ow_sum(w_sum_39_33), .ow_c(w_carry_39_33));
wire w_sum_39_31, w_carry_39_31;
math_adder_carry_save CSA_39_31(.i_a(w_carry_38_45), .i_b(w_carry_38_43), .i_c(w_carry_38_41), .ow_sum(w_sum_39_31), .ow_c(w_carry_39_31));
wire w_sum_39_29, w_carry_39_29;
math_adder_carry_save CSA_39_29(.i_a(w_carry_38_39), .i_b(w_carry_38_37), .i_c(w_carry_38_35), .ow_sum(w_sum_39_29), .ow_c(w_carry_39_29));
wire w_sum_39_27, w_carry_39_27;
math_adder_carry_save CSA_39_27(.i_a(w_carry_38_33), .i_b(w_carry_38_31), .i_c(w_carry_38_29), .ow_sum(w_sum_39_27), .ow_c(w_carry_39_27));
wire w_sum_39_25, w_carry_39_25;
math_adder_carry_save CSA_39_25(.i_a(w_carry_38_27), .i_b(w_carry_38_25), .i_c(w_carry_38_23), .ow_sum(w_sum_39_25), .ow_c(w_carry_39_25));
wire w_sum_39_23, w_carry_39_23;
math_adder_carry_save CSA_39_23(.i_a(w_carry_38_21), .i_b(w_carry_38_19), .i_c(w_carry_38_17), .ow_sum(w_sum_39_23), .ow_c(w_carry_39_23));
wire w_sum_39_21, w_carry_39_21;
math_adder_carry_save CSA_39_21(.i_a(w_carry_38_15), .i_b(w_carry_38_13), .i_c(w_carry_38_11), .ow_sum(w_sum_39_21), .ow_c(w_carry_39_21));
wire w_sum_39_19, w_carry_39_19;
math_adder_carry_save CSA_39_19(.i_a(w_carry_38_9), .i_b(w_carry_38_7), .i_c(w_carry_38_5), .ow_sum(w_sum_39_19), .ow_c(w_carry_39_19));
wire w_sum_39_17, w_carry_39_17;
math_adder_carry_save CSA_39_17(.i_a(w_carry_38_3), .i_b(w_sum_39_49), .i_c(w_sum_39_47), .ow_sum(w_sum_39_17), .ow_c(w_carry_39_17));
wire w_sum_39_15, w_carry_39_15;
math_adder_carry_save CSA_39_15(.i_a(w_sum_39_45), .i_b(w_sum_39_43), .i_c(w_sum_39_41), .ow_sum(w_sum_39_15), .ow_c(w_carry_39_15));
wire w_sum_39_13, w_carry_39_13;
math_adder_carry_save CSA_39_13(.i_a(w_sum_39_39), .i_b(w_sum_39_37), .i_c(w_sum_39_35), .ow_sum(w_sum_39_13), .ow_c(w_carry_39_13));
wire w_sum_39_11, w_carry_39_11;
math_adder_carry_save CSA_39_11(.i_a(w_sum_39_33), .i_b(w_sum_39_31), .i_c(w_sum_39_29), .ow_sum(w_sum_39_11), .ow_c(w_carry_39_11));
wire w_sum_39_9, w_carry_39_9;
math_adder_carry_save CSA_39_9(.i_a(w_sum_39_27), .i_b(w_sum_39_25), .i_c(w_sum_39_23), .ow_sum(w_sum_39_9), .ow_c(w_carry_39_9));
wire w_sum_39_7, w_carry_39_7;
math_adder_carry_save CSA_39_7(.i_a(w_sum_39_21), .i_b(w_sum_39_19), .i_c(w_sum_39_17), .ow_sum(w_sum_39_7), .ow_c(w_carry_39_7));
wire w_sum_39_5, w_carry_39_5;
math_adder_carry_save CSA_39_5(.i_a(w_sum_39_15), .i_b(w_sum_39_13), .i_c(w_sum_39_11), .ow_sum(w_sum_39_5), .ow_c(w_carry_39_5));
wire w_sum_39_3, w_carry_39_3;
math_adder_carry_save CSA_39_3(.i_a(w_sum_39_9), .i_b(w_sum_39_7), .i_c(w_sum_39_5), .ow_sum(w_sum_39_3), .ow_c(w_carry_39_3));
wire w_sum_40_47, w_carry_40_47;
math_adder_carry_save CSA_40_47(.i_a(w_pp_9_31), .i_b(w_pp_10_30), .i_c(w_pp_11_29), .ow_sum(w_sum_40_47), .ow_c(w_carry_40_47));
wire w_sum_40_45, w_carry_40_45;
math_adder_carry_save CSA_40_45(.i_a(w_pp_12_28), .i_b(w_pp_13_27), .i_c(w_pp_14_26), .ow_sum(w_sum_40_45), .ow_c(w_carry_40_45));
wire w_sum_40_43, w_carry_40_43;
math_adder_carry_save CSA_40_43(.i_a(w_pp_15_25), .i_b(w_pp_16_24), .i_c(w_pp_17_23), .ow_sum(w_sum_40_43), .ow_c(w_carry_40_43));
wire w_sum_40_41, w_carry_40_41;
math_adder_carry_save CSA_40_41(.i_a(w_pp_18_22), .i_b(w_pp_19_21), .i_c(w_pp_20_20), .ow_sum(w_sum_40_41), .ow_c(w_carry_40_41));
wire w_sum_40_39, w_carry_40_39;
math_adder_carry_save CSA_40_39(.i_a(w_pp_21_19), .i_b(w_pp_22_18), .i_c(w_pp_23_17), .ow_sum(w_sum_40_39), .ow_c(w_carry_40_39));
wire w_sum_40_37, w_carry_40_37;
math_adder_carry_save CSA_40_37(.i_a(w_pp_24_16), .i_b(w_pp_25_15), .i_c(w_pp_26_14), .ow_sum(w_sum_40_37), .ow_c(w_carry_40_37));
wire w_sum_40_35, w_carry_40_35;
math_adder_carry_save CSA_40_35(.i_a(w_pp_27_13), .i_b(w_pp_28_12), .i_c(w_pp_29_11), .ow_sum(w_sum_40_35), .ow_c(w_carry_40_35));
wire w_sum_40_33, w_carry_40_33;
math_adder_carry_save CSA_40_33(.i_a(w_pp_30_10), .i_b(w_pp_31_9), .i_c(w_carry_39_49), .ow_sum(w_sum_40_33), .ow_c(w_carry_40_33));
wire w_sum_40_31, w_carry_40_31;
math_adder_carry_save CSA_40_31(.i_a(w_carry_39_47), .i_b(w_carry_39_45), .i_c(w_carry_39_43), .ow_sum(w_sum_40_31), .ow_c(w_carry_40_31));
wire w_sum_40_29, w_carry_40_29;
math_adder_carry_save CSA_40_29(.i_a(w_carry_39_41), .i_b(w_carry_39_39), .i_c(w_carry_39_37), .ow_sum(w_sum_40_29), .ow_c(w_carry_40_29));
wire w_sum_40_27, w_carry_40_27;
math_adder_carry_save CSA_40_27(.i_a(w_carry_39_35), .i_b(w_carry_39_33), .i_c(w_carry_39_31), .ow_sum(w_sum_40_27), .ow_c(w_carry_40_27));
wire w_sum_40_25, w_carry_40_25;
math_adder_carry_save CSA_40_25(.i_a(w_carry_39_29), .i_b(w_carry_39_27), .i_c(w_carry_39_25), .ow_sum(w_sum_40_25), .ow_c(w_carry_40_25));
wire w_sum_40_23, w_carry_40_23;
math_adder_carry_save CSA_40_23(.i_a(w_carry_39_23), .i_b(w_carry_39_21), .i_c(w_carry_39_19), .ow_sum(w_sum_40_23), .ow_c(w_carry_40_23));
wire w_sum_40_21, w_carry_40_21;
math_adder_carry_save CSA_40_21(.i_a(w_carry_39_17), .i_b(w_carry_39_15), .i_c(w_carry_39_13), .ow_sum(w_sum_40_21), .ow_c(w_carry_40_21));
wire w_sum_40_19, w_carry_40_19;
math_adder_carry_save CSA_40_19(.i_a(w_carry_39_11), .i_b(w_carry_39_9), .i_c(w_carry_39_7), .ow_sum(w_sum_40_19), .ow_c(w_carry_40_19));
wire w_sum_40_17, w_carry_40_17;
math_adder_carry_save CSA_40_17(.i_a(w_carry_39_5), .i_b(w_carry_39_3), .i_c(w_sum_40_47), .ow_sum(w_sum_40_17), .ow_c(w_carry_40_17));
wire w_sum_40_15, w_carry_40_15;
math_adder_carry_save CSA_40_15(.i_a(w_sum_40_45), .i_b(w_sum_40_43), .i_c(w_sum_40_41), .ow_sum(w_sum_40_15), .ow_c(w_carry_40_15));
wire w_sum_40_13, w_carry_40_13;
math_adder_carry_save CSA_40_13(.i_a(w_sum_40_39), .i_b(w_sum_40_37), .i_c(w_sum_40_35), .ow_sum(w_sum_40_13), .ow_c(w_carry_40_13));
wire w_sum_40_11, w_carry_40_11;
math_adder_carry_save CSA_40_11(.i_a(w_sum_40_33), .i_b(w_sum_40_31), .i_c(w_sum_40_29), .ow_sum(w_sum_40_11), .ow_c(w_carry_40_11));
wire w_sum_40_9, w_carry_40_9;
math_adder_carry_save CSA_40_9(.i_a(w_sum_40_27), .i_b(w_sum_40_25), .i_c(w_sum_40_23), .ow_sum(w_sum_40_9), .ow_c(w_carry_40_9));
wire w_sum_40_7, w_carry_40_7;
math_adder_carry_save CSA_40_7(.i_a(w_sum_40_21), .i_b(w_sum_40_19), .i_c(w_sum_40_17), .ow_sum(w_sum_40_7), .ow_c(w_carry_40_7));
wire w_sum_40_5, w_carry_40_5;
math_adder_carry_save CSA_40_5(.i_a(w_sum_40_15), .i_b(w_sum_40_13), .i_c(w_sum_40_11), .ow_sum(w_sum_40_5), .ow_c(w_carry_40_5));
wire w_sum_40_3, w_carry_40_3;
math_adder_carry_save CSA_40_3(.i_a(w_sum_40_9), .i_b(w_sum_40_7), .i_c(w_sum_40_5), .ow_sum(w_sum_40_3), .ow_c(w_carry_40_3));
wire w_sum_41_45, w_carry_41_45;
math_adder_carry_save CSA_41_45(.i_a(w_pp_10_31), .i_b(w_pp_11_30), .i_c(w_pp_12_29), .ow_sum(w_sum_41_45), .ow_c(w_carry_41_45));
wire w_sum_41_43, w_carry_41_43;
math_adder_carry_save CSA_41_43(.i_a(w_pp_13_28), .i_b(w_pp_14_27), .i_c(w_pp_15_26), .ow_sum(w_sum_41_43), .ow_c(w_carry_41_43));
wire w_sum_41_41, w_carry_41_41;
math_adder_carry_save CSA_41_41(.i_a(w_pp_16_25), .i_b(w_pp_17_24), .i_c(w_pp_18_23), .ow_sum(w_sum_41_41), .ow_c(w_carry_41_41));
wire w_sum_41_39, w_carry_41_39;
math_adder_carry_save CSA_41_39(.i_a(w_pp_19_22), .i_b(w_pp_20_21), .i_c(w_pp_21_20), .ow_sum(w_sum_41_39), .ow_c(w_carry_41_39));
wire w_sum_41_37, w_carry_41_37;
math_adder_carry_save CSA_41_37(.i_a(w_pp_22_19), .i_b(w_pp_23_18), .i_c(w_pp_24_17), .ow_sum(w_sum_41_37), .ow_c(w_carry_41_37));
wire w_sum_41_35, w_carry_41_35;
math_adder_carry_save CSA_41_35(.i_a(w_pp_25_16), .i_b(w_pp_26_15), .i_c(w_pp_27_14), .ow_sum(w_sum_41_35), .ow_c(w_carry_41_35));
wire w_sum_41_33, w_carry_41_33;
math_adder_carry_save CSA_41_33(.i_a(w_pp_28_13), .i_b(w_pp_29_12), .i_c(w_pp_30_11), .ow_sum(w_sum_41_33), .ow_c(w_carry_41_33));
wire w_sum_41_31, w_carry_41_31;
math_adder_carry_save CSA_41_31(.i_a(w_pp_31_10), .i_b(w_carry_40_47), .i_c(w_carry_40_45), .ow_sum(w_sum_41_31), .ow_c(w_carry_41_31));
wire w_sum_41_29, w_carry_41_29;
math_adder_carry_save CSA_41_29(.i_a(w_carry_40_43), .i_b(w_carry_40_41), .i_c(w_carry_40_39), .ow_sum(w_sum_41_29), .ow_c(w_carry_41_29));
wire w_sum_41_27, w_carry_41_27;
math_adder_carry_save CSA_41_27(.i_a(w_carry_40_37), .i_b(w_carry_40_35), .i_c(w_carry_40_33), .ow_sum(w_sum_41_27), .ow_c(w_carry_41_27));
wire w_sum_41_25, w_carry_41_25;
math_adder_carry_save CSA_41_25(.i_a(w_carry_40_31), .i_b(w_carry_40_29), .i_c(w_carry_40_27), .ow_sum(w_sum_41_25), .ow_c(w_carry_41_25));
wire w_sum_41_23, w_carry_41_23;
math_adder_carry_save CSA_41_23(.i_a(w_carry_40_25), .i_b(w_carry_40_23), .i_c(w_carry_40_21), .ow_sum(w_sum_41_23), .ow_c(w_carry_41_23));
wire w_sum_41_21, w_carry_41_21;
math_adder_carry_save CSA_41_21(.i_a(w_carry_40_19), .i_b(w_carry_40_17), .i_c(w_carry_40_15), .ow_sum(w_sum_41_21), .ow_c(w_carry_41_21));
wire w_sum_41_19, w_carry_41_19;
math_adder_carry_save CSA_41_19(.i_a(w_carry_40_13), .i_b(w_carry_40_11), .i_c(w_carry_40_9), .ow_sum(w_sum_41_19), .ow_c(w_carry_41_19));
wire w_sum_41_17, w_carry_41_17;
math_adder_carry_save CSA_41_17(.i_a(w_carry_40_7), .i_b(w_carry_40_5), .i_c(w_carry_40_3), .ow_sum(w_sum_41_17), .ow_c(w_carry_41_17));
wire w_sum_41_15, w_carry_41_15;
math_adder_carry_save CSA_41_15(.i_a(w_sum_41_45), .i_b(w_sum_41_43), .i_c(w_sum_41_41), .ow_sum(w_sum_41_15), .ow_c(w_carry_41_15));
wire w_sum_41_13, w_carry_41_13;
math_adder_carry_save CSA_41_13(.i_a(w_sum_41_39), .i_b(w_sum_41_37), .i_c(w_sum_41_35), .ow_sum(w_sum_41_13), .ow_c(w_carry_41_13));
wire w_sum_41_11, w_carry_41_11;
math_adder_carry_save CSA_41_11(.i_a(w_sum_41_33), .i_b(w_sum_41_31), .i_c(w_sum_41_29), .ow_sum(w_sum_41_11), .ow_c(w_carry_41_11));
wire w_sum_41_9, w_carry_41_9;
math_adder_carry_save CSA_41_9(.i_a(w_sum_41_27), .i_b(w_sum_41_25), .i_c(w_sum_41_23), .ow_sum(w_sum_41_9), .ow_c(w_carry_41_9));
wire w_sum_41_7, w_carry_41_7;
math_adder_carry_save CSA_41_7(.i_a(w_sum_41_21), .i_b(w_sum_41_19), .i_c(w_sum_41_17), .ow_sum(w_sum_41_7), .ow_c(w_carry_41_7));
wire w_sum_41_5, w_carry_41_5;
math_adder_carry_save CSA_41_5(.i_a(w_sum_41_15), .i_b(w_sum_41_13), .i_c(w_sum_41_11), .ow_sum(w_sum_41_5), .ow_c(w_carry_41_5));
wire w_sum_41_3, w_carry_41_3;
math_adder_carry_save CSA_41_3(.i_a(w_sum_41_9), .i_b(w_sum_41_7), .i_c(w_sum_41_5), .ow_sum(w_sum_41_3), .ow_c(w_carry_41_3));
wire w_sum_42_43, w_carry_42_43;
math_adder_carry_save CSA_42_43(.i_a(w_pp_11_31), .i_b(w_pp_12_30), .i_c(w_pp_13_29), .ow_sum(w_sum_42_43), .ow_c(w_carry_42_43));
wire w_sum_42_41, w_carry_42_41;
math_adder_carry_save CSA_42_41(.i_a(w_pp_14_28), .i_b(w_pp_15_27), .i_c(w_pp_16_26), .ow_sum(w_sum_42_41), .ow_c(w_carry_42_41));
wire w_sum_42_39, w_carry_42_39;
math_adder_carry_save CSA_42_39(.i_a(w_pp_17_25), .i_b(w_pp_18_24), .i_c(w_pp_19_23), .ow_sum(w_sum_42_39), .ow_c(w_carry_42_39));
wire w_sum_42_37, w_carry_42_37;
math_adder_carry_save CSA_42_37(.i_a(w_pp_20_22), .i_b(w_pp_21_21), .i_c(w_pp_22_20), .ow_sum(w_sum_42_37), .ow_c(w_carry_42_37));
wire w_sum_42_35, w_carry_42_35;
math_adder_carry_save CSA_42_35(.i_a(w_pp_23_19), .i_b(w_pp_24_18), .i_c(w_pp_25_17), .ow_sum(w_sum_42_35), .ow_c(w_carry_42_35));
wire w_sum_42_33, w_carry_42_33;
math_adder_carry_save CSA_42_33(.i_a(w_pp_26_16), .i_b(w_pp_27_15), .i_c(w_pp_28_14), .ow_sum(w_sum_42_33), .ow_c(w_carry_42_33));
wire w_sum_42_31, w_carry_42_31;
math_adder_carry_save CSA_42_31(.i_a(w_pp_29_13), .i_b(w_pp_30_12), .i_c(w_pp_31_11), .ow_sum(w_sum_42_31), .ow_c(w_carry_42_31));
wire w_sum_42_29, w_carry_42_29;
math_adder_carry_save CSA_42_29(.i_a(w_carry_41_45), .i_b(w_carry_41_43), .i_c(w_carry_41_41), .ow_sum(w_sum_42_29), .ow_c(w_carry_42_29));
wire w_sum_42_27, w_carry_42_27;
math_adder_carry_save CSA_42_27(.i_a(w_carry_41_39), .i_b(w_carry_41_37), .i_c(w_carry_41_35), .ow_sum(w_sum_42_27), .ow_c(w_carry_42_27));
wire w_sum_42_25, w_carry_42_25;
math_adder_carry_save CSA_42_25(.i_a(w_carry_41_33), .i_b(w_carry_41_31), .i_c(w_carry_41_29), .ow_sum(w_sum_42_25), .ow_c(w_carry_42_25));
wire w_sum_42_23, w_carry_42_23;
math_adder_carry_save CSA_42_23(.i_a(w_carry_41_27), .i_b(w_carry_41_25), .i_c(w_carry_41_23), .ow_sum(w_sum_42_23), .ow_c(w_carry_42_23));
wire w_sum_42_21, w_carry_42_21;
math_adder_carry_save CSA_42_21(.i_a(w_carry_41_21), .i_b(w_carry_41_19), .i_c(w_carry_41_17), .ow_sum(w_sum_42_21), .ow_c(w_carry_42_21));
wire w_sum_42_19, w_carry_42_19;
math_adder_carry_save CSA_42_19(.i_a(w_carry_41_15), .i_b(w_carry_41_13), .i_c(w_carry_41_11), .ow_sum(w_sum_42_19), .ow_c(w_carry_42_19));
wire w_sum_42_17, w_carry_42_17;
math_adder_carry_save CSA_42_17(.i_a(w_carry_41_9), .i_b(w_carry_41_7), .i_c(w_carry_41_5), .ow_sum(w_sum_42_17), .ow_c(w_carry_42_17));
wire w_sum_42_15, w_carry_42_15;
math_adder_carry_save CSA_42_15(.i_a(w_carry_41_3), .i_b(w_sum_42_43), .i_c(w_sum_42_41), .ow_sum(w_sum_42_15), .ow_c(w_carry_42_15));
wire w_sum_42_13, w_carry_42_13;
math_adder_carry_save CSA_42_13(.i_a(w_sum_42_39), .i_b(w_sum_42_37), .i_c(w_sum_42_35), .ow_sum(w_sum_42_13), .ow_c(w_carry_42_13));
wire w_sum_42_11, w_carry_42_11;
math_adder_carry_save CSA_42_11(.i_a(w_sum_42_33), .i_b(w_sum_42_31), .i_c(w_sum_42_29), .ow_sum(w_sum_42_11), .ow_c(w_carry_42_11));
wire w_sum_42_9, w_carry_42_9;
math_adder_carry_save CSA_42_9(.i_a(w_sum_42_27), .i_b(w_sum_42_25), .i_c(w_sum_42_23), .ow_sum(w_sum_42_9), .ow_c(w_carry_42_9));
wire w_sum_42_7, w_carry_42_7;
math_adder_carry_save CSA_42_7(.i_a(w_sum_42_21), .i_b(w_sum_42_19), .i_c(w_sum_42_17), .ow_sum(w_sum_42_7), .ow_c(w_carry_42_7));
wire w_sum_42_5, w_carry_42_5;
math_adder_carry_save CSA_42_5(.i_a(w_sum_42_15), .i_b(w_sum_42_13), .i_c(w_sum_42_11), .ow_sum(w_sum_42_5), .ow_c(w_carry_42_5));
wire w_sum_42_3, w_carry_42_3;
math_adder_carry_save CSA_42_3(.i_a(w_sum_42_9), .i_b(w_sum_42_7), .i_c(w_sum_42_5), .ow_sum(w_sum_42_3), .ow_c(w_carry_42_3));
wire w_sum_43_41, w_carry_43_41;
math_adder_carry_save CSA_43_41(.i_a(w_pp_12_31), .i_b(w_pp_13_30), .i_c(w_pp_14_29), .ow_sum(w_sum_43_41), .ow_c(w_carry_43_41));
wire w_sum_43_39, w_carry_43_39;
math_adder_carry_save CSA_43_39(.i_a(w_pp_15_28), .i_b(w_pp_16_27), .i_c(w_pp_17_26), .ow_sum(w_sum_43_39), .ow_c(w_carry_43_39));
wire w_sum_43_37, w_carry_43_37;
math_adder_carry_save CSA_43_37(.i_a(w_pp_18_25), .i_b(w_pp_19_24), .i_c(w_pp_20_23), .ow_sum(w_sum_43_37), .ow_c(w_carry_43_37));
wire w_sum_43_35, w_carry_43_35;
math_adder_carry_save CSA_43_35(.i_a(w_pp_21_22), .i_b(w_pp_22_21), .i_c(w_pp_23_20), .ow_sum(w_sum_43_35), .ow_c(w_carry_43_35));
wire w_sum_43_33, w_carry_43_33;
math_adder_carry_save CSA_43_33(.i_a(w_pp_24_19), .i_b(w_pp_25_18), .i_c(w_pp_26_17), .ow_sum(w_sum_43_33), .ow_c(w_carry_43_33));
wire w_sum_43_31, w_carry_43_31;
math_adder_carry_save CSA_43_31(.i_a(w_pp_27_16), .i_b(w_pp_28_15), .i_c(w_pp_29_14), .ow_sum(w_sum_43_31), .ow_c(w_carry_43_31));
wire w_sum_43_29, w_carry_43_29;
math_adder_carry_save CSA_43_29(.i_a(w_pp_30_13), .i_b(w_pp_31_12), .i_c(w_carry_42_43), .ow_sum(w_sum_43_29), .ow_c(w_carry_43_29));
wire w_sum_43_27, w_carry_43_27;
math_adder_carry_save CSA_43_27(.i_a(w_carry_42_41), .i_b(w_carry_42_39), .i_c(w_carry_42_37), .ow_sum(w_sum_43_27), .ow_c(w_carry_43_27));
wire w_sum_43_25, w_carry_43_25;
math_adder_carry_save CSA_43_25(.i_a(w_carry_42_35), .i_b(w_carry_42_33), .i_c(w_carry_42_31), .ow_sum(w_sum_43_25), .ow_c(w_carry_43_25));
wire w_sum_43_23, w_carry_43_23;
math_adder_carry_save CSA_43_23(.i_a(w_carry_42_29), .i_b(w_carry_42_27), .i_c(w_carry_42_25), .ow_sum(w_sum_43_23), .ow_c(w_carry_43_23));
wire w_sum_43_21, w_carry_43_21;
math_adder_carry_save CSA_43_21(.i_a(w_carry_42_23), .i_b(w_carry_42_21), .i_c(w_carry_42_19), .ow_sum(w_sum_43_21), .ow_c(w_carry_43_21));
wire w_sum_43_19, w_carry_43_19;
math_adder_carry_save CSA_43_19(.i_a(w_carry_42_17), .i_b(w_carry_42_15), .i_c(w_carry_42_13), .ow_sum(w_sum_43_19), .ow_c(w_carry_43_19));
wire w_sum_43_17, w_carry_43_17;
math_adder_carry_save CSA_43_17(.i_a(w_carry_42_11), .i_b(w_carry_42_9), .i_c(w_carry_42_7), .ow_sum(w_sum_43_17), .ow_c(w_carry_43_17));
wire w_sum_43_15, w_carry_43_15;
math_adder_carry_save CSA_43_15(.i_a(w_carry_42_5), .i_b(w_carry_42_3), .i_c(w_sum_43_41), .ow_sum(w_sum_43_15), .ow_c(w_carry_43_15));
wire w_sum_43_13, w_carry_43_13;
math_adder_carry_save CSA_43_13(.i_a(w_sum_43_39), .i_b(w_sum_43_37), .i_c(w_sum_43_35), .ow_sum(w_sum_43_13), .ow_c(w_carry_43_13));
wire w_sum_43_11, w_carry_43_11;
math_adder_carry_save CSA_43_11(.i_a(w_sum_43_33), .i_b(w_sum_43_31), .i_c(w_sum_43_29), .ow_sum(w_sum_43_11), .ow_c(w_carry_43_11));
wire w_sum_43_9, w_carry_43_9;
math_adder_carry_save CSA_43_9(.i_a(w_sum_43_27), .i_b(w_sum_43_25), .i_c(w_sum_43_23), .ow_sum(w_sum_43_9), .ow_c(w_carry_43_9));
wire w_sum_43_7, w_carry_43_7;
math_adder_carry_save CSA_43_7(.i_a(w_sum_43_21), .i_b(w_sum_43_19), .i_c(w_sum_43_17), .ow_sum(w_sum_43_7), .ow_c(w_carry_43_7));
wire w_sum_43_5, w_carry_43_5;
math_adder_carry_save CSA_43_5(.i_a(w_sum_43_15), .i_b(w_sum_43_13), .i_c(w_sum_43_11), .ow_sum(w_sum_43_5), .ow_c(w_carry_43_5));
wire w_sum_43_3, w_carry_43_3;
math_adder_carry_save CSA_43_3(.i_a(w_sum_43_9), .i_b(w_sum_43_7), .i_c(w_sum_43_5), .ow_sum(w_sum_43_3), .ow_c(w_carry_43_3));
wire w_sum_44_39, w_carry_44_39;
math_adder_carry_save CSA_44_39(.i_a(w_pp_13_31), .i_b(w_pp_14_30), .i_c(w_pp_15_29), .ow_sum(w_sum_44_39), .ow_c(w_carry_44_39));
wire w_sum_44_37, w_carry_44_37;
math_adder_carry_save CSA_44_37(.i_a(w_pp_16_28), .i_b(w_pp_17_27), .i_c(w_pp_18_26), .ow_sum(w_sum_44_37), .ow_c(w_carry_44_37));
wire w_sum_44_35, w_carry_44_35;
math_adder_carry_save CSA_44_35(.i_a(w_pp_19_25), .i_b(w_pp_20_24), .i_c(w_pp_21_23), .ow_sum(w_sum_44_35), .ow_c(w_carry_44_35));
wire w_sum_44_33, w_carry_44_33;
math_adder_carry_save CSA_44_33(.i_a(w_pp_22_22), .i_b(w_pp_23_21), .i_c(w_pp_24_20), .ow_sum(w_sum_44_33), .ow_c(w_carry_44_33));
wire w_sum_44_31, w_carry_44_31;
math_adder_carry_save CSA_44_31(.i_a(w_pp_25_19), .i_b(w_pp_26_18), .i_c(w_pp_27_17), .ow_sum(w_sum_44_31), .ow_c(w_carry_44_31));
wire w_sum_44_29, w_carry_44_29;
math_adder_carry_save CSA_44_29(.i_a(w_pp_28_16), .i_b(w_pp_29_15), .i_c(w_pp_30_14), .ow_sum(w_sum_44_29), .ow_c(w_carry_44_29));
wire w_sum_44_27, w_carry_44_27;
math_adder_carry_save CSA_44_27(.i_a(w_pp_31_13), .i_b(w_carry_43_41), .i_c(w_carry_43_39), .ow_sum(w_sum_44_27), .ow_c(w_carry_44_27));
wire w_sum_44_25, w_carry_44_25;
math_adder_carry_save CSA_44_25(.i_a(w_carry_43_37), .i_b(w_carry_43_35), .i_c(w_carry_43_33), .ow_sum(w_sum_44_25), .ow_c(w_carry_44_25));
wire w_sum_44_23, w_carry_44_23;
math_adder_carry_save CSA_44_23(.i_a(w_carry_43_31), .i_b(w_carry_43_29), .i_c(w_carry_43_27), .ow_sum(w_sum_44_23), .ow_c(w_carry_44_23));
wire w_sum_44_21, w_carry_44_21;
math_adder_carry_save CSA_44_21(.i_a(w_carry_43_25), .i_b(w_carry_43_23), .i_c(w_carry_43_21), .ow_sum(w_sum_44_21), .ow_c(w_carry_44_21));
wire w_sum_44_19, w_carry_44_19;
math_adder_carry_save CSA_44_19(.i_a(w_carry_43_19), .i_b(w_carry_43_17), .i_c(w_carry_43_15), .ow_sum(w_sum_44_19), .ow_c(w_carry_44_19));
wire w_sum_44_17, w_carry_44_17;
math_adder_carry_save CSA_44_17(.i_a(w_carry_43_13), .i_b(w_carry_43_11), .i_c(w_carry_43_9), .ow_sum(w_sum_44_17), .ow_c(w_carry_44_17));
wire w_sum_44_15, w_carry_44_15;
math_adder_carry_save CSA_44_15(.i_a(w_carry_43_7), .i_b(w_carry_43_5), .i_c(w_carry_43_3), .ow_sum(w_sum_44_15), .ow_c(w_carry_44_15));
wire w_sum_44_13, w_carry_44_13;
math_adder_carry_save CSA_44_13(.i_a(w_sum_44_39), .i_b(w_sum_44_37), .i_c(w_sum_44_35), .ow_sum(w_sum_44_13), .ow_c(w_carry_44_13));
wire w_sum_44_11, w_carry_44_11;
math_adder_carry_save CSA_44_11(.i_a(w_sum_44_33), .i_b(w_sum_44_31), .i_c(w_sum_44_29), .ow_sum(w_sum_44_11), .ow_c(w_carry_44_11));
wire w_sum_44_9, w_carry_44_9;
math_adder_carry_save CSA_44_9(.i_a(w_sum_44_27), .i_b(w_sum_44_25), .i_c(w_sum_44_23), .ow_sum(w_sum_44_9), .ow_c(w_carry_44_9));
wire w_sum_44_7, w_carry_44_7;
math_adder_carry_save CSA_44_7(.i_a(w_sum_44_21), .i_b(w_sum_44_19), .i_c(w_sum_44_17), .ow_sum(w_sum_44_7), .ow_c(w_carry_44_7));
wire w_sum_44_5, w_carry_44_5;
math_adder_carry_save CSA_44_5(.i_a(w_sum_44_15), .i_b(w_sum_44_13), .i_c(w_sum_44_11), .ow_sum(w_sum_44_5), .ow_c(w_carry_44_5));
wire w_sum_44_3, w_carry_44_3;
math_adder_carry_save CSA_44_3(.i_a(w_sum_44_9), .i_b(w_sum_44_7), .i_c(w_sum_44_5), .ow_sum(w_sum_44_3), .ow_c(w_carry_44_3));
wire w_sum_45_37, w_carry_45_37;
math_adder_carry_save CSA_45_37(.i_a(w_pp_14_31), .i_b(w_pp_15_30), .i_c(w_pp_16_29), .ow_sum(w_sum_45_37), .ow_c(w_carry_45_37));
wire w_sum_45_35, w_carry_45_35;
math_adder_carry_save CSA_45_35(.i_a(w_pp_17_28), .i_b(w_pp_18_27), .i_c(w_pp_19_26), .ow_sum(w_sum_45_35), .ow_c(w_carry_45_35));
wire w_sum_45_33, w_carry_45_33;
math_adder_carry_save CSA_45_33(.i_a(w_pp_20_25), .i_b(w_pp_21_24), .i_c(w_pp_22_23), .ow_sum(w_sum_45_33), .ow_c(w_carry_45_33));
wire w_sum_45_31, w_carry_45_31;
math_adder_carry_save CSA_45_31(.i_a(w_pp_23_22), .i_b(w_pp_24_21), .i_c(w_pp_25_20), .ow_sum(w_sum_45_31), .ow_c(w_carry_45_31));
wire w_sum_45_29, w_carry_45_29;
math_adder_carry_save CSA_45_29(.i_a(w_pp_26_19), .i_b(w_pp_27_18), .i_c(w_pp_28_17), .ow_sum(w_sum_45_29), .ow_c(w_carry_45_29));
wire w_sum_45_27, w_carry_45_27;
math_adder_carry_save CSA_45_27(.i_a(w_pp_29_16), .i_b(w_pp_30_15), .i_c(w_pp_31_14), .ow_sum(w_sum_45_27), .ow_c(w_carry_45_27));
wire w_sum_45_25, w_carry_45_25;
math_adder_carry_save CSA_45_25(.i_a(w_carry_44_39), .i_b(w_carry_44_37), .i_c(w_carry_44_35), .ow_sum(w_sum_45_25), .ow_c(w_carry_45_25));
wire w_sum_45_23, w_carry_45_23;
math_adder_carry_save CSA_45_23(.i_a(w_carry_44_33), .i_b(w_carry_44_31), .i_c(w_carry_44_29), .ow_sum(w_sum_45_23), .ow_c(w_carry_45_23));
wire w_sum_45_21, w_carry_45_21;
math_adder_carry_save CSA_45_21(.i_a(w_carry_44_27), .i_b(w_carry_44_25), .i_c(w_carry_44_23), .ow_sum(w_sum_45_21), .ow_c(w_carry_45_21));
wire w_sum_45_19, w_carry_45_19;
math_adder_carry_save CSA_45_19(.i_a(w_carry_44_21), .i_b(w_carry_44_19), .i_c(w_carry_44_17), .ow_sum(w_sum_45_19), .ow_c(w_carry_45_19));
wire w_sum_45_17, w_carry_45_17;
math_adder_carry_save CSA_45_17(.i_a(w_carry_44_15), .i_b(w_carry_44_13), .i_c(w_carry_44_11), .ow_sum(w_sum_45_17), .ow_c(w_carry_45_17));
wire w_sum_45_15, w_carry_45_15;
math_adder_carry_save CSA_45_15(.i_a(w_carry_44_9), .i_b(w_carry_44_7), .i_c(w_carry_44_5), .ow_sum(w_sum_45_15), .ow_c(w_carry_45_15));
wire w_sum_45_13, w_carry_45_13;
math_adder_carry_save CSA_45_13(.i_a(w_carry_44_3), .i_b(w_sum_45_37), .i_c(w_sum_45_35), .ow_sum(w_sum_45_13), .ow_c(w_carry_45_13));
wire w_sum_45_11, w_carry_45_11;
math_adder_carry_save CSA_45_11(.i_a(w_sum_45_33), .i_b(w_sum_45_31), .i_c(w_sum_45_29), .ow_sum(w_sum_45_11), .ow_c(w_carry_45_11));
wire w_sum_45_9, w_carry_45_9;
math_adder_carry_save CSA_45_9(.i_a(w_sum_45_27), .i_b(w_sum_45_25), .i_c(w_sum_45_23), .ow_sum(w_sum_45_9), .ow_c(w_carry_45_9));
wire w_sum_45_7, w_carry_45_7;
math_adder_carry_save CSA_45_7(.i_a(w_sum_45_21), .i_b(w_sum_45_19), .i_c(w_sum_45_17), .ow_sum(w_sum_45_7), .ow_c(w_carry_45_7));
wire w_sum_45_5, w_carry_45_5;
math_adder_carry_save CSA_45_5(.i_a(w_sum_45_15), .i_b(w_sum_45_13), .i_c(w_sum_45_11), .ow_sum(w_sum_45_5), .ow_c(w_carry_45_5));
wire w_sum_45_3, w_carry_45_3;
math_adder_carry_save CSA_45_3(.i_a(w_sum_45_9), .i_b(w_sum_45_7), .i_c(w_sum_45_5), .ow_sum(w_sum_45_3), .ow_c(w_carry_45_3));
wire w_sum_46_35, w_carry_46_35;
math_adder_carry_save CSA_46_35(.i_a(w_pp_15_31), .i_b(w_pp_16_30), .i_c(w_pp_17_29), .ow_sum(w_sum_46_35), .ow_c(w_carry_46_35));
wire w_sum_46_33, w_carry_46_33;
math_adder_carry_save CSA_46_33(.i_a(w_pp_18_28), .i_b(w_pp_19_27), .i_c(w_pp_20_26), .ow_sum(w_sum_46_33), .ow_c(w_carry_46_33));
wire w_sum_46_31, w_carry_46_31;
math_adder_carry_save CSA_46_31(.i_a(w_pp_21_25), .i_b(w_pp_22_24), .i_c(w_pp_23_23), .ow_sum(w_sum_46_31), .ow_c(w_carry_46_31));
wire w_sum_46_29, w_carry_46_29;
math_adder_carry_save CSA_46_29(.i_a(w_pp_24_22), .i_b(w_pp_25_21), .i_c(w_pp_26_20), .ow_sum(w_sum_46_29), .ow_c(w_carry_46_29));
wire w_sum_46_27, w_carry_46_27;
math_adder_carry_save CSA_46_27(.i_a(w_pp_27_19), .i_b(w_pp_28_18), .i_c(w_pp_29_17), .ow_sum(w_sum_46_27), .ow_c(w_carry_46_27));
wire w_sum_46_25, w_carry_46_25;
math_adder_carry_save CSA_46_25(.i_a(w_pp_30_16), .i_b(w_pp_31_15), .i_c(w_carry_45_37), .ow_sum(w_sum_46_25), .ow_c(w_carry_46_25));
wire w_sum_46_23, w_carry_46_23;
math_adder_carry_save CSA_46_23(.i_a(w_carry_45_35), .i_b(w_carry_45_33), .i_c(w_carry_45_31), .ow_sum(w_sum_46_23), .ow_c(w_carry_46_23));
wire w_sum_46_21, w_carry_46_21;
math_adder_carry_save CSA_46_21(.i_a(w_carry_45_29), .i_b(w_carry_45_27), .i_c(w_carry_45_25), .ow_sum(w_sum_46_21), .ow_c(w_carry_46_21));
wire w_sum_46_19, w_carry_46_19;
math_adder_carry_save CSA_46_19(.i_a(w_carry_45_23), .i_b(w_carry_45_21), .i_c(w_carry_45_19), .ow_sum(w_sum_46_19), .ow_c(w_carry_46_19));
wire w_sum_46_17, w_carry_46_17;
math_adder_carry_save CSA_46_17(.i_a(w_carry_45_17), .i_b(w_carry_45_15), .i_c(w_carry_45_13), .ow_sum(w_sum_46_17), .ow_c(w_carry_46_17));
wire w_sum_46_15, w_carry_46_15;
math_adder_carry_save CSA_46_15(.i_a(w_carry_45_11), .i_b(w_carry_45_9), .i_c(w_carry_45_7), .ow_sum(w_sum_46_15), .ow_c(w_carry_46_15));
wire w_sum_46_13, w_carry_46_13;
math_adder_carry_save CSA_46_13(.i_a(w_carry_45_5), .i_b(w_carry_45_3), .i_c(w_sum_46_35), .ow_sum(w_sum_46_13), .ow_c(w_carry_46_13));
wire w_sum_46_11, w_carry_46_11;
math_adder_carry_save CSA_46_11(.i_a(w_sum_46_33), .i_b(w_sum_46_31), .i_c(w_sum_46_29), .ow_sum(w_sum_46_11), .ow_c(w_carry_46_11));
wire w_sum_46_9, w_carry_46_9;
math_adder_carry_save CSA_46_9(.i_a(w_sum_46_27), .i_b(w_sum_46_25), .i_c(w_sum_46_23), .ow_sum(w_sum_46_9), .ow_c(w_carry_46_9));
wire w_sum_46_7, w_carry_46_7;
math_adder_carry_save CSA_46_7(.i_a(w_sum_46_21), .i_b(w_sum_46_19), .i_c(w_sum_46_17), .ow_sum(w_sum_46_7), .ow_c(w_carry_46_7));
wire w_sum_46_5, w_carry_46_5;
math_adder_carry_save CSA_46_5(.i_a(w_sum_46_15), .i_b(w_sum_46_13), .i_c(w_sum_46_11), .ow_sum(w_sum_46_5), .ow_c(w_carry_46_5));
wire w_sum_46_3, w_carry_46_3;
math_adder_carry_save CSA_46_3(.i_a(w_sum_46_9), .i_b(w_sum_46_7), .i_c(w_sum_46_5), .ow_sum(w_sum_46_3), .ow_c(w_carry_46_3));
wire w_sum_47_33, w_carry_47_33;
math_adder_carry_save CSA_47_33(.i_a(w_pp_16_31), .i_b(w_pp_17_30), .i_c(w_pp_18_29), .ow_sum(w_sum_47_33), .ow_c(w_carry_47_33));
wire w_sum_47_31, w_carry_47_31;
math_adder_carry_save CSA_47_31(.i_a(w_pp_19_28), .i_b(w_pp_20_27), .i_c(w_pp_21_26), .ow_sum(w_sum_47_31), .ow_c(w_carry_47_31));
wire w_sum_47_29, w_carry_47_29;
math_adder_carry_save CSA_47_29(.i_a(w_pp_22_25), .i_b(w_pp_23_24), .i_c(w_pp_24_23), .ow_sum(w_sum_47_29), .ow_c(w_carry_47_29));
wire w_sum_47_27, w_carry_47_27;
math_adder_carry_save CSA_47_27(.i_a(w_pp_25_22), .i_b(w_pp_26_21), .i_c(w_pp_27_20), .ow_sum(w_sum_47_27), .ow_c(w_carry_47_27));
wire w_sum_47_25, w_carry_47_25;
math_adder_carry_save CSA_47_25(.i_a(w_pp_28_19), .i_b(w_pp_29_18), .i_c(w_pp_30_17), .ow_sum(w_sum_47_25), .ow_c(w_carry_47_25));
wire w_sum_47_23, w_carry_47_23;
math_adder_carry_save CSA_47_23(.i_a(w_pp_31_16), .i_b(w_carry_46_35), .i_c(w_carry_46_33), .ow_sum(w_sum_47_23), .ow_c(w_carry_47_23));
wire w_sum_47_21, w_carry_47_21;
math_adder_carry_save CSA_47_21(.i_a(w_carry_46_31), .i_b(w_carry_46_29), .i_c(w_carry_46_27), .ow_sum(w_sum_47_21), .ow_c(w_carry_47_21));
wire w_sum_47_19, w_carry_47_19;
math_adder_carry_save CSA_47_19(.i_a(w_carry_46_25), .i_b(w_carry_46_23), .i_c(w_carry_46_21), .ow_sum(w_sum_47_19), .ow_c(w_carry_47_19));
wire w_sum_47_17, w_carry_47_17;
math_adder_carry_save CSA_47_17(.i_a(w_carry_46_19), .i_b(w_carry_46_17), .i_c(w_carry_46_15), .ow_sum(w_sum_47_17), .ow_c(w_carry_47_17));
wire w_sum_47_15, w_carry_47_15;
math_adder_carry_save CSA_47_15(.i_a(w_carry_46_13), .i_b(w_carry_46_11), .i_c(w_carry_46_9), .ow_sum(w_sum_47_15), .ow_c(w_carry_47_15));
wire w_sum_47_13, w_carry_47_13;
math_adder_carry_save CSA_47_13(.i_a(w_carry_46_7), .i_b(w_carry_46_5), .i_c(w_carry_46_3), .ow_sum(w_sum_47_13), .ow_c(w_carry_47_13));
wire w_sum_47_11, w_carry_47_11;
math_adder_carry_save CSA_47_11(.i_a(w_sum_47_33), .i_b(w_sum_47_31), .i_c(w_sum_47_29), .ow_sum(w_sum_47_11), .ow_c(w_carry_47_11));
wire w_sum_47_9, w_carry_47_9;
math_adder_carry_save CSA_47_9(.i_a(w_sum_47_27), .i_b(w_sum_47_25), .i_c(w_sum_47_23), .ow_sum(w_sum_47_9), .ow_c(w_carry_47_9));
wire w_sum_47_7, w_carry_47_7;
math_adder_carry_save CSA_47_7(.i_a(w_sum_47_21), .i_b(w_sum_47_19), .i_c(w_sum_47_17), .ow_sum(w_sum_47_7), .ow_c(w_carry_47_7));
wire w_sum_47_5, w_carry_47_5;
math_adder_carry_save CSA_47_5(.i_a(w_sum_47_15), .i_b(w_sum_47_13), .i_c(w_sum_47_11), .ow_sum(w_sum_47_5), .ow_c(w_carry_47_5));
wire w_sum_47_3, w_carry_47_3;
math_adder_carry_save CSA_47_3(.i_a(w_sum_47_9), .i_b(w_sum_47_7), .i_c(w_sum_47_5), .ow_sum(w_sum_47_3), .ow_c(w_carry_47_3));
wire w_sum_48_31, w_carry_48_31;
math_adder_carry_save CSA_48_31(.i_a(w_pp_17_31), .i_b(w_pp_18_30), .i_c(w_pp_19_29), .ow_sum(w_sum_48_31), .ow_c(w_carry_48_31));
wire w_sum_48_29, w_carry_48_29;
math_adder_carry_save CSA_48_29(.i_a(w_pp_20_28), .i_b(w_pp_21_27), .i_c(w_pp_22_26), .ow_sum(w_sum_48_29), .ow_c(w_carry_48_29));
wire w_sum_48_27, w_carry_48_27;
math_adder_carry_save CSA_48_27(.i_a(w_pp_23_25), .i_b(w_pp_24_24), .i_c(w_pp_25_23), .ow_sum(w_sum_48_27), .ow_c(w_carry_48_27));
wire w_sum_48_25, w_carry_48_25;
math_adder_carry_save CSA_48_25(.i_a(w_pp_26_22), .i_b(w_pp_27_21), .i_c(w_pp_28_20), .ow_sum(w_sum_48_25), .ow_c(w_carry_48_25));
wire w_sum_48_23, w_carry_48_23;
math_adder_carry_save CSA_48_23(.i_a(w_pp_29_19), .i_b(w_pp_30_18), .i_c(w_pp_31_17), .ow_sum(w_sum_48_23), .ow_c(w_carry_48_23));
wire w_sum_48_21, w_carry_48_21;
math_adder_carry_save CSA_48_21(.i_a(w_carry_47_33), .i_b(w_carry_47_31), .i_c(w_carry_47_29), .ow_sum(w_sum_48_21), .ow_c(w_carry_48_21));
wire w_sum_48_19, w_carry_48_19;
math_adder_carry_save CSA_48_19(.i_a(w_carry_47_27), .i_b(w_carry_47_25), .i_c(w_carry_47_23), .ow_sum(w_sum_48_19), .ow_c(w_carry_48_19));
wire w_sum_48_17, w_carry_48_17;
math_adder_carry_save CSA_48_17(.i_a(w_carry_47_21), .i_b(w_carry_47_19), .i_c(w_carry_47_17), .ow_sum(w_sum_48_17), .ow_c(w_carry_48_17));
wire w_sum_48_15, w_carry_48_15;
math_adder_carry_save CSA_48_15(.i_a(w_carry_47_15), .i_b(w_carry_47_13), .i_c(w_carry_47_11), .ow_sum(w_sum_48_15), .ow_c(w_carry_48_15));
wire w_sum_48_13, w_carry_48_13;
math_adder_carry_save CSA_48_13(.i_a(w_carry_47_9), .i_b(w_carry_47_7), .i_c(w_carry_47_5), .ow_sum(w_sum_48_13), .ow_c(w_carry_48_13));
wire w_sum_48_11, w_carry_48_11;
math_adder_carry_save CSA_48_11(.i_a(w_carry_47_3), .i_b(w_sum_48_31), .i_c(w_sum_48_29), .ow_sum(w_sum_48_11), .ow_c(w_carry_48_11));
wire w_sum_48_9, w_carry_48_9;
math_adder_carry_save CSA_48_9(.i_a(w_sum_48_27), .i_b(w_sum_48_25), .i_c(w_sum_48_23), .ow_sum(w_sum_48_9), .ow_c(w_carry_48_9));
wire w_sum_48_7, w_carry_48_7;
math_adder_carry_save CSA_48_7(.i_a(w_sum_48_21), .i_b(w_sum_48_19), .i_c(w_sum_48_17), .ow_sum(w_sum_48_7), .ow_c(w_carry_48_7));
wire w_sum_48_5, w_carry_48_5;
math_adder_carry_save CSA_48_5(.i_a(w_sum_48_15), .i_b(w_sum_48_13), .i_c(w_sum_48_11), .ow_sum(w_sum_48_5), .ow_c(w_carry_48_5));
wire w_sum_48_3, w_carry_48_3;
math_adder_carry_save CSA_48_3(.i_a(w_sum_48_9), .i_b(w_sum_48_7), .i_c(w_sum_48_5), .ow_sum(w_sum_48_3), .ow_c(w_carry_48_3));
wire w_sum_49_29, w_carry_49_29;
math_adder_carry_save CSA_49_29(.i_a(w_pp_18_31), .i_b(w_pp_19_30), .i_c(w_pp_20_29), .ow_sum(w_sum_49_29), .ow_c(w_carry_49_29));
wire w_sum_49_27, w_carry_49_27;
math_adder_carry_save CSA_49_27(.i_a(w_pp_21_28), .i_b(w_pp_22_27), .i_c(w_pp_23_26), .ow_sum(w_sum_49_27), .ow_c(w_carry_49_27));
wire w_sum_49_25, w_carry_49_25;
math_adder_carry_save CSA_49_25(.i_a(w_pp_24_25), .i_b(w_pp_25_24), .i_c(w_pp_26_23), .ow_sum(w_sum_49_25), .ow_c(w_carry_49_25));
wire w_sum_49_23, w_carry_49_23;
math_adder_carry_save CSA_49_23(.i_a(w_pp_27_22), .i_b(w_pp_28_21), .i_c(w_pp_29_20), .ow_sum(w_sum_49_23), .ow_c(w_carry_49_23));
wire w_sum_49_21, w_carry_49_21;
math_adder_carry_save CSA_49_21(.i_a(w_pp_30_19), .i_b(w_pp_31_18), .i_c(w_carry_48_31), .ow_sum(w_sum_49_21), .ow_c(w_carry_49_21));
wire w_sum_49_19, w_carry_49_19;
math_adder_carry_save CSA_49_19(.i_a(w_carry_48_29), .i_b(w_carry_48_27), .i_c(w_carry_48_25), .ow_sum(w_sum_49_19), .ow_c(w_carry_49_19));
wire w_sum_49_17, w_carry_49_17;
math_adder_carry_save CSA_49_17(.i_a(w_carry_48_23), .i_b(w_carry_48_21), .i_c(w_carry_48_19), .ow_sum(w_sum_49_17), .ow_c(w_carry_49_17));
wire w_sum_49_15, w_carry_49_15;
math_adder_carry_save CSA_49_15(.i_a(w_carry_48_17), .i_b(w_carry_48_15), .i_c(w_carry_48_13), .ow_sum(w_sum_49_15), .ow_c(w_carry_49_15));
wire w_sum_49_13, w_carry_49_13;
math_adder_carry_save CSA_49_13(.i_a(w_carry_48_11), .i_b(w_carry_48_9), .i_c(w_carry_48_7), .ow_sum(w_sum_49_13), .ow_c(w_carry_49_13));
wire w_sum_49_11, w_carry_49_11;
math_adder_carry_save CSA_49_11(.i_a(w_carry_48_5), .i_b(w_carry_48_3), .i_c(w_sum_49_29), .ow_sum(w_sum_49_11), .ow_c(w_carry_49_11));
wire w_sum_49_9, w_carry_49_9;
math_adder_carry_save CSA_49_9(.i_a(w_sum_49_27), .i_b(w_sum_49_25), .i_c(w_sum_49_23), .ow_sum(w_sum_49_9), .ow_c(w_carry_49_9));
wire w_sum_49_7, w_carry_49_7;
math_adder_carry_save CSA_49_7(.i_a(w_sum_49_21), .i_b(w_sum_49_19), .i_c(w_sum_49_17), .ow_sum(w_sum_49_7), .ow_c(w_carry_49_7));
wire w_sum_49_5, w_carry_49_5;
math_adder_carry_save CSA_49_5(.i_a(w_sum_49_15), .i_b(w_sum_49_13), .i_c(w_sum_49_11), .ow_sum(w_sum_49_5), .ow_c(w_carry_49_5));
wire w_sum_49_3, w_carry_49_3;
math_adder_carry_save CSA_49_3(.i_a(w_sum_49_9), .i_b(w_sum_49_7), .i_c(w_sum_49_5), .ow_sum(w_sum_49_3), .ow_c(w_carry_49_3));
wire w_sum_50_27, w_carry_50_27;
math_adder_carry_save CSA_50_27(.i_a(w_pp_19_31), .i_b(w_pp_20_30), .i_c(w_pp_21_29), .ow_sum(w_sum_50_27), .ow_c(w_carry_50_27));
wire w_sum_50_25, w_carry_50_25;
math_adder_carry_save CSA_50_25(.i_a(w_pp_22_28), .i_b(w_pp_23_27), .i_c(w_pp_24_26), .ow_sum(w_sum_50_25), .ow_c(w_carry_50_25));
wire w_sum_50_23, w_carry_50_23;
math_adder_carry_save CSA_50_23(.i_a(w_pp_25_25), .i_b(w_pp_26_24), .i_c(w_pp_27_23), .ow_sum(w_sum_50_23), .ow_c(w_carry_50_23));
wire w_sum_50_21, w_carry_50_21;
math_adder_carry_save CSA_50_21(.i_a(w_pp_28_22), .i_b(w_pp_29_21), .i_c(w_pp_30_20), .ow_sum(w_sum_50_21), .ow_c(w_carry_50_21));
wire w_sum_50_19, w_carry_50_19;
math_adder_carry_save CSA_50_19(.i_a(w_pp_31_19), .i_b(w_carry_49_29), .i_c(w_carry_49_27), .ow_sum(w_sum_50_19), .ow_c(w_carry_50_19));
wire w_sum_50_17, w_carry_50_17;
math_adder_carry_save CSA_50_17(.i_a(w_carry_49_25), .i_b(w_carry_49_23), .i_c(w_carry_49_21), .ow_sum(w_sum_50_17), .ow_c(w_carry_50_17));
wire w_sum_50_15, w_carry_50_15;
math_adder_carry_save CSA_50_15(.i_a(w_carry_49_19), .i_b(w_carry_49_17), .i_c(w_carry_49_15), .ow_sum(w_sum_50_15), .ow_c(w_carry_50_15));
wire w_sum_50_13, w_carry_50_13;
math_adder_carry_save CSA_50_13(.i_a(w_carry_49_13), .i_b(w_carry_49_11), .i_c(w_carry_49_9), .ow_sum(w_sum_50_13), .ow_c(w_carry_50_13));
wire w_sum_50_11, w_carry_50_11;
math_adder_carry_save CSA_50_11(.i_a(w_carry_49_7), .i_b(w_carry_49_5), .i_c(w_carry_49_3), .ow_sum(w_sum_50_11), .ow_c(w_carry_50_11));
wire w_sum_50_9, w_carry_50_9;
math_adder_carry_save CSA_50_9(.i_a(w_sum_50_27), .i_b(w_sum_50_25), .i_c(w_sum_50_23), .ow_sum(w_sum_50_9), .ow_c(w_carry_50_9));
wire w_sum_50_7, w_carry_50_7;
math_adder_carry_save CSA_50_7(.i_a(w_sum_50_21), .i_b(w_sum_50_19), .i_c(w_sum_50_17), .ow_sum(w_sum_50_7), .ow_c(w_carry_50_7));
wire w_sum_50_5, w_carry_50_5;
math_adder_carry_save CSA_50_5(.i_a(w_sum_50_15), .i_b(w_sum_50_13), .i_c(w_sum_50_11), .ow_sum(w_sum_50_5), .ow_c(w_carry_50_5));
wire w_sum_50_3, w_carry_50_3;
math_adder_carry_save CSA_50_3(.i_a(w_sum_50_9), .i_b(w_sum_50_7), .i_c(w_sum_50_5), .ow_sum(w_sum_50_3), .ow_c(w_carry_50_3));
wire w_sum_51_25, w_carry_51_25;
math_adder_carry_save CSA_51_25(.i_a(w_pp_20_31), .i_b(w_pp_21_30), .i_c(w_pp_22_29), .ow_sum(w_sum_51_25), .ow_c(w_carry_51_25));
wire w_sum_51_23, w_carry_51_23;
math_adder_carry_save CSA_51_23(.i_a(w_pp_23_28), .i_b(w_pp_24_27), .i_c(w_pp_25_26), .ow_sum(w_sum_51_23), .ow_c(w_carry_51_23));
wire w_sum_51_21, w_carry_51_21;
math_adder_carry_save CSA_51_21(.i_a(w_pp_26_25), .i_b(w_pp_27_24), .i_c(w_pp_28_23), .ow_sum(w_sum_51_21), .ow_c(w_carry_51_21));
wire w_sum_51_19, w_carry_51_19;
math_adder_carry_save CSA_51_19(.i_a(w_pp_29_22), .i_b(w_pp_30_21), .i_c(w_pp_31_20), .ow_sum(w_sum_51_19), .ow_c(w_carry_51_19));
wire w_sum_51_17, w_carry_51_17;
math_adder_carry_save CSA_51_17(.i_a(w_carry_50_27), .i_b(w_carry_50_25), .i_c(w_carry_50_23), .ow_sum(w_sum_51_17), .ow_c(w_carry_51_17));
wire w_sum_51_15, w_carry_51_15;
math_adder_carry_save CSA_51_15(.i_a(w_carry_50_21), .i_b(w_carry_50_19), .i_c(w_carry_50_17), .ow_sum(w_sum_51_15), .ow_c(w_carry_51_15));
wire w_sum_51_13, w_carry_51_13;
math_adder_carry_save CSA_51_13(.i_a(w_carry_50_15), .i_b(w_carry_50_13), .i_c(w_carry_50_11), .ow_sum(w_sum_51_13), .ow_c(w_carry_51_13));
wire w_sum_51_11, w_carry_51_11;
math_adder_carry_save CSA_51_11(.i_a(w_carry_50_9), .i_b(w_carry_50_7), .i_c(w_carry_50_5), .ow_sum(w_sum_51_11), .ow_c(w_carry_51_11));
wire w_sum_51_9, w_carry_51_9;
math_adder_carry_save CSA_51_9(.i_a(w_carry_50_3), .i_b(w_sum_51_25), .i_c(w_sum_51_23), .ow_sum(w_sum_51_9), .ow_c(w_carry_51_9));
wire w_sum_51_7, w_carry_51_7;
math_adder_carry_save CSA_51_7(.i_a(w_sum_51_21), .i_b(w_sum_51_19), .i_c(w_sum_51_17), .ow_sum(w_sum_51_7), .ow_c(w_carry_51_7));
wire w_sum_51_5, w_carry_51_5;
math_adder_carry_save CSA_51_5(.i_a(w_sum_51_15), .i_b(w_sum_51_13), .i_c(w_sum_51_11), .ow_sum(w_sum_51_5), .ow_c(w_carry_51_5));
wire w_sum_51_3, w_carry_51_3;
math_adder_carry_save CSA_51_3(.i_a(w_sum_51_9), .i_b(w_sum_51_7), .i_c(w_sum_51_5), .ow_sum(w_sum_51_3), .ow_c(w_carry_51_3));
wire w_sum_52_23, w_carry_52_23;
math_adder_carry_save CSA_52_23(.i_a(w_pp_21_31), .i_b(w_pp_22_30), .i_c(w_pp_23_29), .ow_sum(w_sum_52_23), .ow_c(w_carry_52_23));
wire w_sum_52_21, w_carry_52_21;
math_adder_carry_save CSA_52_21(.i_a(w_pp_24_28), .i_b(w_pp_25_27), .i_c(w_pp_26_26), .ow_sum(w_sum_52_21), .ow_c(w_carry_52_21));
wire w_sum_52_19, w_carry_52_19;
math_adder_carry_save CSA_52_19(.i_a(w_pp_27_25), .i_b(w_pp_28_24), .i_c(w_pp_29_23), .ow_sum(w_sum_52_19), .ow_c(w_carry_52_19));
wire w_sum_52_17, w_carry_52_17;
math_adder_carry_save CSA_52_17(.i_a(w_pp_30_22), .i_b(w_pp_31_21), .i_c(w_carry_51_25), .ow_sum(w_sum_52_17), .ow_c(w_carry_52_17));
wire w_sum_52_15, w_carry_52_15;
math_adder_carry_save CSA_52_15(.i_a(w_carry_51_23), .i_b(w_carry_51_21), .i_c(w_carry_51_19), .ow_sum(w_sum_52_15), .ow_c(w_carry_52_15));
wire w_sum_52_13, w_carry_52_13;
math_adder_carry_save CSA_52_13(.i_a(w_carry_51_17), .i_b(w_carry_51_15), .i_c(w_carry_51_13), .ow_sum(w_sum_52_13), .ow_c(w_carry_52_13));
wire w_sum_52_11, w_carry_52_11;
math_adder_carry_save CSA_52_11(.i_a(w_carry_51_11), .i_b(w_carry_51_9), .i_c(w_carry_51_7), .ow_sum(w_sum_52_11), .ow_c(w_carry_52_11));
wire w_sum_52_9, w_carry_52_9;
math_adder_carry_save CSA_52_9(.i_a(w_carry_51_5), .i_b(w_carry_51_3), .i_c(w_sum_52_23), .ow_sum(w_sum_52_9), .ow_c(w_carry_52_9));
wire w_sum_52_7, w_carry_52_7;
math_adder_carry_save CSA_52_7(.i_a(w_sum_52_21), .i_b(w_sum_52_19), .i_c(w_sum_52_17), .ow_sum(w_sum_52_7), .ow_c(w_carry_52_7));
wire w_sum_52_5, w_carry_52_5;
math_adder_carry_save CSA_52_5(.i_a(w_sum_52_15), .i_b(w_sum_52_13), .i_c(w_sum_52_11), .ow_sum(w_sum_52_5), .ow_c(w_carry_52_5));
wire w_sum_52_3, w_carry_52_3;
math_adder_carry_save CSA_52_3(.i_a(w_sum_52_9), .i_b(w_sum_52_7), .i_c(w_sum_52_5), .ow_sum(w_sum_52_3), .ow_c(w_carry_52_3));
wire w_sum_53_21, w_carry_53_21;
math_adder_carry_save CSA_53_21(.i_a(w_pp_22_31), .i_b(w_pp_23_30), .i_c(w_pp_24_29), .ow_sum(w_sum_53_21), .ow_c(w_carry_53_21));
wire w_sum_53_19, w_carry_53_19;
math_adder_carry_save CSA_53_19(.i_a(w_pp_25_28), .i_b(w_pp_26_27), .i_c(w_pp_27_26), .ow_sum(w_sum_53_19), .ow_c(w_carry_53_19));
wire w_sum_53_17, w_carry_53_17;
math_adder_carry_save CSA_53_17(.i_a(w_pp_28_25), .i_b(w_pp_29_24), .i_c(w_pp_30_23), .ow_sum(w_sum_53_17), .ow_c(w_carry_53_17));
wire w_sum_53_15, w_carry_53_15;
math_adder_carry_save CSA_53_15(.i_a(w_pp_31_22), .i_b(w_carry_52_23), .i_c(w_carry_52_21), .ow_sum(w_sum_53_15), .ow_c(w_carry_53_15));
wire w_sum_53_13, w_carry_53_13;
math_adder_carry_save CSA_53_13(.i_a(w_carry_52_19), .i_b(w_carry_52_17), .i_c(w_carry_52_15), .ow_sum(w_sum_53_13), .ow_c(w_carry_53_13));
wire w_sum_53_11, w_carry_53_11;
math_adder_carry_save CSA_53_11(.i_a(w_carry_52_13), .i_b(w_carry_52_11), .i_c(w_carry_52_9), .ow_sum(w_sum_53_11), .ow_c(w_carry_53_11));
wire w_sum_53_9, w_carry_53_9;
math_adder_carry_save CSA_53_9(.i_a(w_carry_52_7), .i_b(w_carry_52_5), .i_c(w_carry_52_3), .ow_sum(w_sum_53_9), .ow_c(w_carry_53_9));
wire w_sum_53_7, w_carry_53_7;
math_adder_carry_save CSA_53_7(.i_a(w_sum_53_21), .i_b(w_sum_53_19), .i_c(w_sum_53_17), .ow_sum(w_sum_53_7), .ow_c(w_carry_53_7));
wire w_sum_53_5, w_carry_53_5;
math_adder_carry_save CSA_53_5(.i_a(w_sum_53_15), .i_b(w_sum_53_13), .i_c(w_sum_53_11), .ow_sum(w_sum_53_5), .ow_c(w_carry_53_5));
wire w_sum_53_3, w_carry_53_3;
math_adder_carry_save CSA_53_3(.i_a(w_sum_53_9), .i_b(w_sum_53_7), .i_c(w_sum_53_5), .ow_sum(w_sum_53_3), .ow_c(w_carry_53_3));
wire w_sum_54_19, w_carry_54_19;
math_adder_carry_save CSA_54_19(.i_a(w_pp_23_31), .i_b(w_pp_24_30), .i_c(w_pp_25_29), .ow_sum(w_sum_54_19), .ow_c(w_carry_54_19));
wire w_sum_54_17, w_carry_54_17;
math_adder_carry_save CSA_54_17(.i_a(w_pp_26_28), .i_b(w_pp_27_27), .i_c(w_pp_28_26), .ow_sum(w_sum_54_17), .ow_c(w_carry_54_17));
wire w_sum_54_15, w_carry_54_15;
math_adder_carry_save CSA_54_15(.i_a(w_pp_29_25), .i_b(w_pp_30_24), .i_c(w_pp_31_23), .ow_sum(w_sum_54_15), .ow_c(w_carry_54_15));
wire w_sum_54_13, w_carry_54_13;
math_adder_carry_save CSA_54_13(.i_a(w_carry_53_21), .i_b(w_carry_53_19), .i_c(w_carry_53_17), .ow_sum(w_sum_54_13), .ow_c(w_carry_54_13));
wire w_sum_54_11, w_carry_54_11;
math_adder_carry_save CSA_54_11(.i_a(w_carry_53_15), .i_b(w_carry_53_13), .i_c(w_carry_53_11), .ow_sum(w_sum_54_11), .ow_c(w_carry_54_11));
wire w_sum_54_9, w_carry_54_9;
math_adder_carry_save CSA_54_9(.i_a(w_carry_53_9), .i_b(w_carry_53_7), .i_c(w_carry_53_5), .ow_sum(w_sum_54_9), .ow_c(w_carry_54_9));
wire w_sum_54_7, w_carry_54_7;
math_adder_carry_save CSA_54_7(.i_a(w_carry_53_3), .i_b(w_sum_54_19), .i_c(w_sum_54_17), .ow_sum(w_sum_54_7), .ow_c(w_carry_54_7));
wire w_sum_54_5, w_carry_54_5;
math_adder_carry_save CSA_54_5(.i_a(w_sum_54_15), .i_b(w_sum_54_13), .i_c(w_sum_54_11), .ow_sum(w_sum_54_5), .ow_c(w_carry_54_5));
wire w_sum_54_3, w_carry_54_3;
math_adder_carry_save CSA_54_3(.i_a(w_sum_54_9), .i_b(w_sum_54_7), .i_c(w_sum_54_5), .ow_sum(w_sum_54_3), .ow_c(w_carry_54_3));
wire w_sum_55_17, w_carry_55_17;
math_adder_carry_save CSA_55_17(.i_a(w_pp_24_31), .i_b(w_pp_25_30), .i_c(w_pp_26_29), .ow_sum(w_sum_55_17), .ow_c(w_carry_55_17));
wire w_sum_55_15, w_carry_55_15;
math_adder_carry_save CSA_55_15(.i_a(w_pp_27_28), .i_b(w_pp_28_27), .i_c(w_pp_29_26), .ow_sum(w_sum_55_15), .ow_c(w_carry_55_15));
wire w_sum_55_13, w_carry_55_13;
math_adder_carry_save CSA_55_13(.i_a(w_pp_30_25), .i_b(w_pp_31_24), .i_c(w_carry_54_19), .ow_sum(w_sum_55_13), .ow_c(w_carry_55_13));
wire w_sum_55_11, w_carry_55_11;
math_adder_carry_save CSA_55_11(.i_a(w_carry_54_17), .i_b(w_carry_54_15), .i_c(w_carry_54_13), .ow_sum(w_sum_55_11), .ow_c(w_carry_55_11));
wire w_sum_55_9, w_carry_55_9;
math_adder_carry_save CSA_55_9(.i_a(w_carry_54_11), .i_b(w_carry_54_9), .i_c(w_carry_54_7), .ow_sum(w_sum_55_9), .ow_c(w_carry_55_9));
wire w_sum_55_7, w_carry_55_7;
math_adder_carry_save CSA_55_7(.i_a(w_carry_54_5), .i_b(w_carry_54_3), .i_c(w_sum_55_17), .ow_sum(w_sum_55_7), .ow_c(w_carry_55_7));
wire w_sum_55_5, w_carry_55_5;
math_adder_carry_save CSA_55_5(.i_a(w_sum_55_15), .i_b(w_sum_55_13), .i_c(w_sum_55_11), .ow_sum(w_sum_55_5), .ow_c(w_carry_55_5));
wire w_sum_55_3, w_carry_55_3;
math_adder_carry_save CSA_55_3(.i_a(w_sum_55_9), .i_b(w_sum_55_7), .i_c(w_sum_55_5), .ow_sum(w_sum_55_3), .ow_c(w_carry_55_3));
wire w_sum_56_15, w_carry_56_15;
math_adder_carry_save CSA_56_15(.i_a(w_pp_25_31), .i_b(w_pp_26_30), .i_c(w_pp_27_29), .ow_sum(w_sum_56_15), .ow_c(w_carry_56_15));
wire w_sum_56_13, w_carry_56_13;
math_adder_carry_save CSA_56_13(.i_a(w_pp_28_28), .i_b(w_pp_29_27), .i_c(w_pp_30_26), .ow_sum(w_sum_56_13), .ow_c(w_carry_56_13));
wire w_sum_56_11, w_carry_56_11;
math_adder_carry_save CSA_56_11(.i_a(w_pp_31_25), .i_b(w_carry_55_17), .i_c(w_carry_55_15), .ow_sum(w_sum_56_11), .ow_c(w_carry_56_11));
wire w_sum_56_9, w_carry_56_9;
math_adder_carry_save CSA_56_9(.i_a(w_carry_55_13), .i_b(w_carry_55_11), .i_c(w_carry_55_9), .ow_sum(w_sum_56_9), .ow_c(w_carry_56_9));
wire w_sum_56_7, w_carry_56_7;
math_adder_carry_save CSA_56_7(.i_a(w_carry_55_7), .i_b(w_carry_55_5), .i_c(w_carry_55_3), .ow_sum(w_sum_56_7), .ow_c(w_carry_56_7));
wire w_sum_56_5, w_carry_56_5;
math_adder_carry_save CSA_56_5(.i_a(w_sum_56_15), .i_b(w_sum_56_13), .i_c(w_sum_56_11), .ow_sum(w_sum_56_5), .ow_c(w_carry_56_5));
wire w_sum_56_3, w_carry_56_3;
math_adder_carry_save CSA_56_3(.i_a(w_sum_56_9), .i_b(w_sum_56_7), .i_c(w_sum_56_5), .ow_sum(w_sum_56_3), .ow_c(w_carry_56_3));
wire w_sum_57_13, w_carry_57_13;
math_adder_carry_save CSA_57_13(.i_a(w_pp_26_31), .i_b(w_pp_27_30), .i_c(w_pp_28_29), .ow_sum(w_sum_57_13), .ow_c(w_carry_57_13));
wire w_sum_57_11, w_carry_57_11;
math_adder_carry_save CSA_57_11(.i_a(w_pp_29_28), .i_b(w_pp_30_27), .i_c(w_pp_31_26), .ow_sum(w_sum_57_11), .ow_c(w_carry_57_11));
wire w_sum_57_9, w_carry_57_9;
math_adder_carry_save CSA_57_9(.i_a(w_carry_56_15), .i_b(w_carry_56_13), .i_c(w_carry_56_11), .ow_sum(w_sum_57_9), .ow_c(w_carry_57_9));
wire w_sum_57_7, w_carry_57_7;
math_adder_carry_save CSA_57_7(.i_a(w_carry_56_9), .i_b(w_carry_56_7), .i_c(w_carry_56_5), .ow_sum(w_sum_57_7), .ow_c(w_carry_57_7));
wire w_sum_57_5, w_carry_57_5;
math_adder_carry_save CSA_57_5(.i_a(w_carry_56_3), .i_b(w_sum_57_13), .i_c(w_sum_57_11), .ow_sum(w_sum_57_5), .ow_c(w_carry_57_5));
wire w_sum_57_3, w_carry_57_3;
math_adder_carry_save CSA_57_3(.i_a(w_sum_57_9), .i_b(w_sum_57_7), .i_c(w_sum_57_5), .ow_sum(w_sum_57_3), .ow_c(w_carry_57_3));
wire w_sum_58_11, w_carry_58_11;
math_adder_carry_save CSA_58_11(.i_a(w_pp_27_31), .i_b(w_pp_28_30), .i_c(w_pp_29_29), .ow_sum(w_sum_58_11), .ow_c(w_carry_58_11));
wire w_sum_58_9, w_carry_58_9;
math_adder_carry_save CSA_58_9(.i_a(w_pp_30_28), .i_b(w_pp_31_27), .i_c(w_carry_57_13), .ow_sum(w_sum_58_9), .ow_c(w_carry_58_9));
wire w_sum_58_7, w_carry_58_7;
math_adder_carry_save CSA_58_7(.i_a(w_carry_57_11), .i_b(w_carry_57_9), .i_c(w_carry_57_7), .ow_sum(w_sum_58_7), .ow_c(w_carry_58_7));
wire w_sum_58_5, w_carry_58_5;
math_adder_carry_save CSA_58_5(.i_a(w_carry_57_5), .i_b(w_carry_57_3), .i_c(w_sum_58_11), .ow_sum(w_sum_58_5), .ow_c(w_carry_58_5));
wire w_sum_58_3, w_carry_58_3;
math_adder_carry_save CSA_58_3(.i_a(w_sum_58_9), .i_b(w_sum_58_7), .i_c(w_sum_58_5), .ow_sum(w_sum_58_3), .ow_c(w_carry_58_3));
wire w_sum_59_9, w_carry_59_9;
math_adder_carry_save CSA_59_9(.i_a(w_pp_28_31), .i_b(w_pp_29_30), .i_c(w_pp_30_29), .ow_sum(w_sum_59_9), .ow_c(w_carry_59_9));
wire w_sum_59_7, w_carry_59_7;
math_adder_carry_save CSA_59_7(.i_a(w_pp_31_28), .i_b(w_carry_58_11), .i_c(w_carry_58_9), .ow_sum(w_sum_59_7), .ow_c(w_carry_59_7));
wire w_sum_59_5, w_carry_59_5;
math_adder_carry_save CSA_59_5(.i_a(w_carry_58_7), .i_b(w_carry_58_5), .i_c(w_carry_58_3), .ow_sum(w_sum_59_5), .ow_c(w_carry_59_5));
wire w_sum_59_3, w_carry_59_3;
math_adder_carry_save CSA_59_3(.i_a(w_sum_59_9), .i_b(w_sum_59_7), .i_c(w_sum_59_5), .ow_sum(w_sum_59_3), .ow_c(w_carry_59_3));
wire w_sum_60_7, w_carry_60_7;
math_adder_carry_save CSA_60_7(.i_a(w_pp_29_31), .i_b(w_pp_30_30), .i_c(w_pp_31_29), .ow_sum(w_sum_60_7), .ow_c(w_carry_60_7));
wire w_sum_60_5, w_carry_60_5;
math_adder_carry_save CSA_60_5(.i_a(w_carry_59_9), .i_b(w_carry_59_7), .i_c(w_carry_59_5), .ow_sum(w_sum_60_5), .ow_c(w_carry_60_5));
wire w_sum_60_3, w_carry_60_3;
math_adder_carry_save CSA_60_3(.i_a(w_carry_59_3), .i_b(w_sum_60_7), .i_c(w_sum_60_5), .ow_sum(w_sum_60_3), .ow_c(w_carry_60_3));
wire w_sum_61_5, w_carry_61_5;
math_adder_carry_save CSA_61_5(.i_a(w_pp_30_31), .i_b(w_pp_31_30), .i_c(w_carry_60_7), .ow_sum(w_sum_61_5), .ow_c(w_carry_61_5));
wire w_sum_61_3, w_carry_61_3;
math_adder_carry_save CSA_61_3(.i_a(w_carry_60_5), .i_b(w_carry_60_3), .i_c(w_sum_61_5), .ow_sum(w_sum_61_3), .ow_c(w_carry_61_3));
wire w_sum_62_3, w_carry_62_3;
math_adder_carry_save CSA_62_3(.i_a(w_pp_31_31), .i_b(w_carry_61_5), .i_c(w_carry_61_3), .ow_sum(w_sum_62_3), .ow_c(w_carry_62_3));

// Final product assignment
assign ow_product[0] = w_pp_0_0;
assign ow_product[1] = w_sum_1_2;
assign ow_product[2] = w_sum_2_2;
assign ow_product[3] = w_sum_3_2;
assign ow_product[4] = w_sum_4_2;
assign ow_product[5] = w_sum_5_2;
assign ow_product[6] = w_sum_6_2;
assign ow_product[7] = w_sum_7_2;
assign ow_product[8] = w_sum_8_2;
assign ow_product[9] = w_sum_9_2;
assign ow_product[10] = w_sum_10_2;
assign ow_product[11] = w_sum_11_2;
assign ow_product[12] = w_sum_12_2;
assign ow_product[13] = w_sum_13_2;
assign ow_product[14] = w_sum_14_2;
assign ow_product[15] = w_sum_15_2;
assign ow_product[16] = w_sum_16_2;
assign ow_product[17] = w_sum_17_2;
assign ow_product[18] = w_sum_18_2;
assign ow_product[19] = w_sum_19_2;
assign ow_product[20] = w_sum_20_2;
assign ow_product[21] = w_sum_21_2;
assign ow_product[22] = w_sum_22_2;
assign ow_product[23] = w_sum_23_2;
assign ow_product[24] = w_sum_24_2;
assign ow_product[25] = w_sum_25_2;
assign ow_product[26] = w_sum_26_2;
assign ow_product[27] = w_sum_27_2;
assign ow_product[28] = w_sum_28_2;
assign ow_product[29] = w_sum_29_2;
assign ow_product[30] = w_sum_30_2;
assign ow_product[31] = w_sum_31_2;
assign ow_product[32] = w_sum_32_2;
assign ow_product[33] = w_sum_33_3;
assign ow_product[34] = w_sum_34_3;
assign ow_product[35] = w_sum_35_3;
assign ow_product[36] = w_sum_36_3;
assign ow_product[37] = w_sum_37_3;
assign ow_product[38] = w_sum_38_3;
assign ow_product[39] = w_sum_39_3;
assign ow_product[40] = w_sum_40_3;
assign ow_product[41] = w_sum_41_3;
assign ow_product[42] = w_sum_42_3;
assign ow_product[43] = w_sum_43_3;
assign ow_product[44] = w_sum_44_3;
assign ow_product[45] = w_sum_45_3;
assign ow_product[46] = w_sum_46_3;
assign ow_product[47] = w_sum_47_3;
assign ow_product[48] = w_sum_48_3;
assign ow_product[49] = w_sum_49_3;
assign ow_product[50] = w_sum_50_3;
assign ow_product[51] = w_sum_51_3;
assign ow_product[52] = w_sum_52_3;
assign ow_product[53] = w_sum_53_3;
assign ow_product[54] = w_sum_54_3;
assign ow_product[55] = w_sum_55_3;
assign ow_product[56] = w_sum_56_3;
assign ow_product[57] = w_sum_57_3;
assign ow_product[58] = w_sum_58_3;
assign ow_product[59] = w_sum_59_3;
assign ow_product[60] = w_sum_60_3;
assign ow_product[61] = w_sum_61_3;
assign ow_product[62] = w_sum_62_3;
assign ow_product[63] = w_carry_62_3;


    // Debug purposes
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_wallace_tree_csa_32);
    end
                
endmodule : math_multiplier_wallace_tree_csa_32
