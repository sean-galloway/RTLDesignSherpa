//      // verilator_coverage annotation
        // SPDX-License-Identifier: MIT
        // SPDX-FileCopyrightText: 2024-2025 sean galloway
        //
        // RTL Design Sherpa - Industry-Standard RTL Design and Verification
        // https://github.com/sean-galloway/RTLDesignSherpa
        //
        // Module: math_addsub_full_nbit
        // Purpose: Math Addsub Full Nbit module
        //
        // Documentation: rtl/common/PRD.md
        // Subsystem: common
        //
        // Author: sean galloway
        // Created: 2025-10-18
        
        `timescale 1ns / 1ps
        
        module math_addsub_full_nbit #(
            parameter int N = 4
        ) (
%000001     input  logic [N-1:0] i_a,
 000031     input  logic [N-1:0] i_b,
 000511     input  logic         i_c,      // 0 for add, 1 for subtract
 000240     output logic [N-1:0] ow_sum,
 000241     output logic         ow_carry  // Final carry-out
        );
        
 000223     logic [  N:0] w_c;  // array for internal carries
 000256     logic [N-1:0] w_ip;  // array XORing i_c and i_b
        
            genvar i;
            generate
                for (i = 0; i < N; i++) begin : gen_xor
                    assign w_ip[i] = i_b[i] ^ i_c;
                end
            endgenerate
        
            assign w_c[0] = i_c;
        
            generate
                for (i = 0; i < N; i++) begin : gen_full_adders
                    math_adder_full fa (
                        .i_a     (i_a[i]),
                        .i_b     (w_ip[i]),
                        .i_c     (w_c[i]),
                        .ow_sum  (ow_sum[i]),
                        .ow_carry(w_c[i+1])
                    );
                end
            endgenerate
        
            assign ow_carry = w_c[N];  // output the final carry or borrow
        
        endmodule : math_addsub_full_nbit
        
