`timescale 1ns / 1ps

module math_multiplier_dadda_tree_016 (
    input  [15:0] i_multiplier,
    input  [15:0] i_multiplicand,
    output [31:0] ow_product
);

// Partial products generation
wire w_pp_00_00 = i_multiplier[ 0] & i_multiplicand[ 0];
wire w_pp_00_01 = i_multiplier[ 0] & i_multiplicand[ 1];
wire w_pp_00_02 = i_multiplier[ 0] & i_multiplicand[ 2];
wire w_pp_00_03 = i_multiplier[ 0] & i_multiplicand[ 3];
wire w_pp_00_04 = i_multiplier[ 0] & i_multiplicand[ 4];
wire w_pp_00_05 = i_multiplier[ 0] & i_multiplicand[ 5];
wire w_pp_00_06 = i_multiplier[ 0] & i_multiplicand[ 6];
wire w_pp_00_07 = i_multiplier[ 0] & i_multiplicand[ 7];
wire w_pp_00_08 = i_multiplier[ 0] & i_multiplicand[ 8];
wire w_pp_00_09 = i_multiplier[ 0] & i_multiplicand[ 9];
wire w_pp_00_10 = i_multiplier[ 0] & i_multiplicand[10];
wire w_pp_00_11 = i_multiplier[ 0] & i_multiplicand[11];
wire w_pp_00_12 = i_multiplier[ 0] & i_multiplicand[12];
wire w_pp_00_13 = i_multiplier[ 0] & i_multiplicand[13];
wire w_pp_00_14 = i_multiplier[ 0] & i_multiplicand[14];
wire w_pp_00_15 = i_multiplier[ 0] & i_multiplicand[15];
wire w_pp_01_00 = i_multiplier[ 1] & i_multiplicand[ 0];
wire w_pp_01_01 = i_multiplier[ 1] & i_multiplicand[ 1];
wire w_pp_01_02 = i_multiplier[ 1] & i_multiplicand[ 2];
wire w_pp_01_03 = i_multiplier[ 1] & i_multiplicand[ 3];
wire w_pp_01_04 = i_multiplier[ 1] & i_multiplicand[ 4];
wire w_pp_01_05 = i_multiplier[ 1] & i_multiplicand[ 5];
wire w_pp_01_06 = i_multiplier[ 1] & i_multiplicand[ 6];
wire w_pp_01_07 = i_multiplier[ 1] & i_multiplicand[ 7];
wire w_pp_01_08 = i_multiplier[ 1] & i_multiplicand[ 8];
wire w_pp_01_09 = i_multiplier[ 1] & i_multiplicand[ 9];
wire w_pp_01_10 = i_multiplier[ 1] & i_multiplicand[10];
wire w_pp_01_11 = i_multiplier[ 1] & i_multiplicand[11];
wire w_pp_01_12 = i_multiplier[ 1] & i_multiplicand[12];
wire w_pp_01_13 = i_multiplier[ 1] & i_multiplicand[13];
wire w_pp_01_14 = i_multiplier[ 1] & i_multiplicand[14];
wire w_pp_01_15 = i_multiplier[ 1] & i_multiplicand[15];
wire w_pp_02_00 = i_multiplier[ 2] & i_multiplicand[ 0];
wire w_pp_02_01 = i_multiplier[ 2] & i_multiplicand[ 1];
wire w_pp_02_02 = i_multiplier[ 2] & i_multiplicand[ 2];
wire w_pp_02_03 = i_multiplier[ 2] & i_multiplicand[ 3];
wire w_pp_02_04 = i_multiplier[ 2] & i_multiplicand[ 4];
wire w_pp_02_05 = i_multiplier[ 2] & i_multiplicand[ 5];
wire w_pp_02_06 = i_multiplier[ 2] & i_multiplicand[ 6];
wire w_pp_02_07 = i_multiplier[ 2] & i_multiplicand[ 7];
wire w_pp_02_08 = i_multiplier[ 2] & i_multiplicand[ 8];
wire w_pp_02_09 = i_multiplier[ 2] & i_multiplicand[ 9];
wire w_pp_02_10 = i_multiplier[ 2] & i_multiplicand[10];
wire w_pp_02_11 = i_multiplier[ 2] & i_multiplicand[11];
wire w_pp_02_12 = i_multiplier[ 2] & i_multiplicand[12];
wire w_pp_02_13 = i_multiplier[ 2] & i_multiplicand[13];
wire w_pp_02_14 = i_multiplier[ 2] & i_multiplicand[14];
wire w_pp_02_15 = i_multiplier[ 2] & i_multiplicand[15];
wire w_pp_03_00 = i_multiplier[ 3] & i_multiplicand[ 0];
wire w_pp_03_01 = i_multiplier[ 3] & i_multiplicand[ 1];
wire w_pp_03_02 = i_multiplier[ 3] & i_multiplicand[ 2];
wire w_pp_03_03 = i_multiplier[ 3] & i_multiplicand[ 3];
wire w_pp_03_04 = i_multiplier[ 3] & i_multiplicand[ 4];
wire w_pp_03_05 = i_multiplier[ 3] & i_multiplicand[ 5];
wire w_pp_03_06 = i_multiplier[ 3] & i_multiplicand[ 6];
wire w_pp_03_07 = i_multiplier[ 3] & i_multiplicand[ 7];
wire w_pp_03_08 = i_multiplier[ 3] & i_multiplicand[ 8];
wire w_pp_03_09 = i_multiplier[ 3] & i_multiplicand[ 9];
wire w_pp_03_10 = i_multiplier[ 3] & i_multiplicand[10];
wire w_pp_03_11 = i_multiplier[ 3] & i_multiplicand[11];
wire w_pp_03_12 = i_multiplier[ 3] & i_multiplicand[12];
wire w_pp_03_13 = i_multiplier[ 3] & i_multiplicand[13];
wire w_pp_03_14 = i_multiplier[ 3] & i_multiplicand[14];
wire w_pp_03_15 = i_multiplier[ 3] & i_multiplicand[15];
wire w_pp_04_00 = i_multiplier[ 4] & i_multiplicand[ 0];
wire w_pp_04_01 = i_multiplier[ 4] & i_multiplicand[ 1];
wire w_pp_04_02 = i_multiplier[ 4] & i_multiplicand[ 2];
wire w_pp_04_03 = i_multiplier[ 4] & i_multiplicand[ 3];
wire w_pp_04_04 = i_multiplier[ 4] & i_multiplicand[ 4];
wire w_pp_04_05 = i_multiplier[ 4] & i_multiplicand[ 5];
wire w_pp_04_06 = i_multiplier[ 4] & i_multiplicand[ 6];
wire w_pp_04_07 = i_multiplier[ 4] & i_multiplicand[ 7];
wire w_pp_04_08 = i_multiplier[ 4] & i_multiplicand[ 8];
wire w_pp_04_09 = i_multiplier[ 4] & i_multiplicand[ 9];
wire w_pp_04_10 = i_multiplier[ 4] & i_multiplicand[10];
wire w_pp_04_11 = i_multiplier[ 4] & i_multiplicand[11];
wire w_pp_04_12 = i_multiplier[ 4] & i_multiplicand[12];
wire w_pp_04_13 = i_multiplier[ 4] & i_multiplicand[13];
wire w_pp_04_14 = i_multiplier[ 4] & i_multiplicand[14];
wire w_pp_04_15 = i_multiplier[ 4] & i_multiplicand[15];
wire w_pp_05_00 = i_multiplier[ 5] & i_multiplicand[ 0];
wire w_pp_05_01 = i_multiplier[ 5] & i_multiplicand[ 1];
wire w_pp_05_02 = i_multiplier[ 5] & i_multiplicand[ 2];
wire w_pp_05_03 = i_multiplier[ 5] & i_multiplicand[ 3];
wire w_pp_05_04 = i_multiplier[ 5] & i_multiplicand[ 4];
wire w_pp_05_05 = i_multiplier[ 5] & i_multiplicand[ 5];
wire w_pp_05_06 = i_multiplier[ 5] & i_multiplicand[ 6];
wire w_pp_05_07 = i_multiplier[ 5] & i_multiplicand[ 7];
wire w_pp_05_08 = i_multiplier[ 5] & i_multiplicand[ 8];
wire w_pp_05_09 = i_multiplier[ 5] & i_multiplicand[ 9];
wire w_pp_05_10 = i_multiplier[ 5] & i_multiplicand[10];
wire w_pp_05_11 = i_multiplier[ 5] & i_multiplicand[11];
wire w_pp_05_12 = i_multiplier[ 5] & i_multiplicand[12];
wire w_pp_05_13 = i_multiplier[ 5] & i_multiplicand[13];
wire w_pp_05_14 = i_multiplier[ 5] & i_multiplicand[14];
wire w_pp_05_15 = i_multiplier[ 5] & i_multiplicand[15];
wire w_pp_06_00 = i_multiplier[ 6] & i_multiplicand[ 0];
wire w_pp_06_01 = i_multiplier[ 6] & i_multiplicand[ 1];
wire w_pp_06_02 = i_multiplier[ 6] & i_multiplicand[ 2];
wire w_pp_06_03 = i_multiplier[ 6] & i_multiplicand[ 3];
wire w_pp_06_04 = i_multiplier[ 6] & i_multiplicand[ 4];
wire w_pp_06_05 = i_multiplier[ 6] & i_multiplicand[ 5];
wire w_pp_06_06 = i_multiplier[ 6] & i_multiplicand[ 6];
wire w_pp_06_07 = i_multiplier[ 6] & i_multiplicand[ 7];
wire w_pp_06_08 = i_multiplier[ 6] & i_multiplicand[ 8];
wire w_pp_06_09 = i_multiplier[ 6] & i_multiplicand[ 9];
wire w_pp_06_10 = i_multiplier[ 6] & i_multiplicand[10];
wire w_pp_06_11 = i_multiplier[ 6] & i_multiplicand[11];
wire w_pp_06_12 = i_multiplier[ 6] & i_multiplicand[12];
wire w_pp_06_13 = i_multiplier[ 6] & i_multiplicand[13];
wire w_pp_06_14 = i_multiplier[ 6] & i_multiplicand[14];
wire w_pp_06_15 = i_multiplier[ 6] & i_multiplicand[15];
wire w_pp_07_00 = i_multiplier[ 7] & i_multiplicand[ 0];
wire w_pp_07_01 = i_multiplier[ 7] & i_multiplicand[ 1];
wire w_pp_07_02 = i_multiplier[ 7] & i_multiplicand[ 2];
wire w_pp_07_03 = i_multiplier[ 7] & i_multiplicand[ 3];
wire w_pp_07_04 = i_multiplier[ 7] & i_multiplicand[ 4];
wire w_pp_07_05 = i_multiplier[ 7] & i_multiplicand[ 5];
wire w_pp_07_06 = i_multiplier[ 7] & i_multiplicand[ 6];
wire w_pp_07_07 = i_multiplier[ 7] & i_multiplicand[ 7];
wire w_pp_07_08 = i_multiplier[ 7] & i_multiplicand[ 8];
wire w_pp_07_09 = i_multiplier[ 7] & i_multiplicand[ 9];
wire w_pp_07_10 = i_multiplier[ 7] & i_multiplicand[10];
wire w_pp_07_11 = i_multiplier[ 7] & i_multiplicand[11];
wire w_pp_07_12 = i_multiplier[ 7] & i_multiplicand[12];
wire w_pp_07_13 = i_multiplier[ 7] & i_multiplicand[13];
wire w_pp_07_14 = i_multiplier[ 7] & i_multiplicand[14];
wire w_pp_07_15 = i_multiplier[ 7] & i_multiplicand[15];
wire w_pp_08_00 = i_multiplier[ 8] & i_multiplicand[ 0];
wire w_pp_08_01 = i_multiplier[ 8] & i_multiplicand[ 1];
wire w_pp_08_02 = i_multiplier[ 8] & i_multiplicand[ 2];
wire w_pp_08_03 = i_multiplier[ 8] & i_multiplicand[ 3];
wire w_pp_08_04 = i_multiplier[ 8] & i_multiplicand[ 4];
wire w_pp_08_05 = i_multiplier[ 8] & i_multiplicand[ 5];
wire w_pp_08_06 = i_multiplier[ 8] & i_multiplicand[ 6];
wire w_pp_08_07 = i_multiplier[ 8] & i_multiplicand[ 7];
wire w_pp_08_08 = i_multiplier[ 8] & i_multiplicand[ 8];
wire w_pp_08_09 = i_multiplier[ 8] & i_multiplicand[ 9];
wire w_pp_08_10 = i_multiplier[ 8] & i_multiplicand[10];
wire w_pp_08_11 = i_multiplier[ 8] & i_multiplicand[11];
wire w_pp_08_12 = i_multiplier[ 8] & i_multiplicand[12];
wire w_pp_08_13 = i_multiplier[ 8] & i_multiplicand[13];
wire w_pp_08_14 = i_multiplier[ 8] & i_multiplicand[14];
wire w_pp_08_15 = i_multiplier[ 8] & i_multiplicand[15];
wire w_pp_09_00 = i_multiplier[ 9] & i_multiplicand[ 0];
wire w_pp_09_01 = i_multiplier[ 9] & i_multiplicand[ 1];
wire w_pp_09_02 = i_multiplier[ 9] & i_multiplicand[ 2];
wire w_pp_09_03 = i_multiplier[ 9] & i_multiplicand[ 3];
wire w_pp_09_04 = i_multiplier[ 9] & i_multiplicand[ 4];
wire w_pp_09_05 = i_multiplier[ 9] & i_multiplicand[ 5];
wire w_pp_09_06 = i_multiplier[ 9] & i_multiplicand[ 6];
wire w_pp_09_07 = i_multiplier[ 9] & i_multiplicand[ 7];
wire w_pp_09_08 = i_multiplier[ 9] & i_multiplicand[ 8];
wire w_pp_09_09 = i_multiplier[ 9] & i_multiplicand[ 9];
wire w_pp_09_10 = i_multiplier[ 9] & i_multiplicand[10];
wire w_pp_09_11 = i_multiplier[ 9] & i_multiplicand[11];
wire w_pp_09_12 = i_multiplier[ 9] & i_multiplicand[12];
wire w_pp_09_13 = i_multiplier[ 9] & i_multiplicand[13];
wire w_pp_09_14 = i_multiplier[ 9] & i_multiplicand[14];
wire w_pp_09_15 = i_multiplier[ 9] & i_multiplicand[15];
wire w_pp_10_00 = i_multiplier[10] & i_multiplicand[ 0];
wire w_pp_10_01 = i_multiplier[10] & i_multiplicand[ 1];
wire w_pp_10_02 = i_multiplier[10] & i_multiplicand[ 2];
wire w_pp_10_03 = i_multiplier[10] & i_multiplicand[ 3];
wire w_pp_10_04 = i_multiplier[10] & i_multiplicand[ 4];
wire w_pp_10_05 = i_multiplier[10] & i_multiplicand[ 5];
wire w_pp_10_06 = i_multiplier[10] & i_multiplicand[ 6];
wire w_pp_10_07 = i_multiplier[10] & i_multiplicand[ 7];
wire w_pp_10_08 = i_multiplier[10] & i_multiplicand[ 8];
wire w_pp_10_09 = i_multiplier[10] & i_multiplicand[ 9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_11_00 = i_multiplier[11] & i_multiplicand[ 0];
wire w_pp_11_01 = i_multiplier[11] & i_multiplicand[ 1];
wire w_pp_11_02 = i_multiplier[11] & i_multiplicand[ 2];
wire w_pp_11_03 = i_multiplier[11] & i_multiplicand[ 3];
wire w_pp_11_04 = i_multiplier[11] & i_multiplicand[ 4];
wire w_pp_11_05 = i_multiplier[11] & i_multiplicand[ 5];
wire w_pp_11_06 = i_multiplier[11] & i_multiplicand[ 6];
wire w_pp_11_07 = i_multiplier[11] & i_multiplicand[ 7];
wire w_pp_11_08 = i_multiplier[11] & i_multiplicand[ 8];
wire w_pp_11_09 = i_multiplier[11] & i_multiplicand[ 9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_12_00 = i_multiplier[12] & i_multiplicand[ 0];
wire w_pp_12_01 = i_multiplier[12] & i_multiplicand[ 1];
wire w_pp_12_02 = i_multiplier[12] & i_multiplicand[ 2];
wire w_pp_12_03 = i_multiplier[12] & i_multiplicand[ 3];
wire w_pp_12_04 = i_multiplier[12] & i_multiplicand[ 4];
wire w_pp_12_05 = i_multiplier[12] & i_multiplicand[ 5];
wire w_pp_12_06 = i_multiplier[12] & i_multiplicand[ 6];
wire w_pp_12_07 = i_multiplier[12] & i_multiplicand[ 7];
wire w_pp_12_08 = i_multiplier[12] & i_multiplicand[ 8];
wire w_pp_12_09 = i_multiplier[12] & i_multiplicand[ 9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_13_00 = i_multiplier[13] & i_multiplicand[ 0];
wire w_pp_13_01 = i_multiplier[13] & i_multiplicand[ 1];
wire w_pp_13_02 = i_multiplier[13] & i_multiplicand[ 2];
wire w_pp_13_03 = i_multiplier[13] & i_multiplicand[ 3];
wire w_pp_13_04 = i_multiplier[13] & i_multiplicand[ 4];
wire w_pp_13_05 = i_multiplier[13] & i_multiplicand[ 5];
wire w_pp_13_06 = i_multiplier[13] & i_multiplicand[ 6];
wire w_pp_13_07 = i_multiplier[13] & i_multiplicand[ 7];
wire w_pp_13_08 = i_multiplier[13] & i_multiplicand[ 8];
wire w_pp_13_09 = i_multiplier[13] & i_multiplicand[ 9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_14_00 = i_multiplier[14] & i_multiplicand[ 0];
wire w_pp_14_01 = i_multiplier[14] & i_multiplicand[ 1];
wire w_pp_14_02 = i_multiplier[14] & i_multiplicand[ 2];
wire w_pp_14_03 = i_multiplier[14] & i_multiplicand[ 3];
wire w_pp_14_04 = i_multiplier[14] & i_multiplicand[ 4];
wire w_pp_14_05 = i_multiplier[14] & i_multiplicand[ 5];
wire w_pp_14_06 = i_multiplier[14] & i_multiplicand[ 6];
wire w_pp_14_07 = i_multiplier[14] & i_multiplicand[ 7];
wire w_pp_14_08 = i_multiplier[14] & i_multiplicand[ 8];
wire w_pp_14_09 = i_multiplier[14] & i_multiplicand[ 9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_15_00 = i_multiplier[15] & i_multiplicand[ 0];
wire w_pp_15_01 = i_multiplier[15] & i_multiplicand[ 1];
wire w_pp_15_02 = i_multiplier[15] & i_multiplicand[ 2];
wire w_pp_15_03 = i_multiplier[15] & i_multiplicand[ 3];
wire w_pp_15_04 = i_multiplier[15] & i_multiplicand[ 4];
wire w_pp_15_05 = i_multiplier[15] & i_multiplicand[ 5];
wire w_pp_15_06 = i_multiplier[15] & i_multiplicand[ 6];
wire w_pp_15_07 = i_multiplier[15] & i_multiplicand[ 7];
wire w_pp_15_08 = i_multiplier[15] & i_multiplicand[ 8];
wire w_pp_15_09 = i_multiplier[15] & i_multiplicand[ 9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];

// Stage: 0, Max Height: 12
wire w_sum_0, w_carry_0;
math_adder_half HA_0(.i_a(w_pp_00_12), .i_b(w_pp_01_11), .ow_sum(w_sum_0), .ow_carry(w_carry_0));
wire w_sum_1, w_carry_1;
math_adder_carry_save CSA_1(.i_a(w_pp_00_13), .i_b(w_pp_01_12), .i_c(w_pp_02_11), .ow_sum(w_sum_1), .ow_carry(w_carry_1));
wire w_sum_2, w_carry_2;
math_adder_half HA_2(.i_a(w_pp_03_10), .i_b(w_pp_04_09), .ow_sum(w_sum_2), .ow_carry(w_carry_2));
wire w_sum_3, w_carry_3;
math_adder_carry_save CSA_3(.i_a(w_pp_00_14), .i_b(w_pp_01_13), .i_c(w_pp_02_12), .ow_sum(w_sum_3), .ow_carry(w_carry_3));
wire w_sum_4, w_carry_4;
math_adder_carry_save CSA_4(.i_a(w_pp_03_11), .i_b(w_pp_04_10), .i_c(w_pp_05_09), .ow_sum(w_sum_4), .ow_carry(w_carry_4));
wire w_sum_5, w_carry_5;
math_adder_half HA_5(.i_a(w_pp_06_08), .i_b(w_pp_07_07), .ow_sum(w_sum_5), .ow_carry(w_carry_5));
wire w_sum_6, w_carry_6;
math_adder_carry_save CSA_6(.i_a(w_pp_00_15), .i_b(w_pp_01_14), .i_c(w_pp_02_13), .ow_sum(w_sum_6), .ow_carry(w_carry_6));
wire w_sum_7, w_carry_7;
math_adder_carry_save CSA_7(.i_a(w_pp_03_12), .i_b(w_pp_04_11), .i_c(w_pp_05_10), .ow_sum(w_sum_7), .ow_carry(w_carry_7));
wire w_sum_8, w_carry_8;
math_adder_carry_save CSA_8(.i_a(w_pp_06_09), .i_b(w_pp_07_08), .i_c(w_pp_08_07), .ow_sum(w_sum_8), .ow_carry(w_carry_8));
wire w_sum_9, w_carry_9;
math_adder_half HA_9(.i_a(w_pp_09_06), .i_b(w_pp_10_05), .ow_sum(w_sum_9), .ow_carry(w_carry_9));
wire w_sum_10, w_carry_10;
math_adder_carry_save CSA_10(.i_a(w_pp_01_15), .i_b(w_pp_02_14), .i_c(w_pp_03_13), .ow_sum(w_sum_10), .ow_carry(w_carry_10));
wire w_sum_11, w_carry_11;
math_adder_carry_save CSA_11(.i_a(w_pp_04_12), .i_b(w_pp_05_11), .i_c(w_pp_06_10), .ow_sum(w_sum_11), .ow_carry(w_carry_11));
wire w_sum_12, w_carry_12;
math_adder_carry_save CSA_12(.i_a(w_pp_07_09), .i_b(w_pp_08_08), .i_c(w_pp_09_07), .ow_sum(w_sum_12), .ow_carry(w_carry_12));
wire w_sum_13, w_carry_13;
math_adder_half HA_13(.i_a(w_pp_10_06), .i_b(w_pp_11_05), .ow_sum(w_sum_13), .ow_carry(w_carry_13));
wire w_sum_14, w_carry_14;
math_adder_carry_save CSA_14(.i_a(w_pp_02_15), .i_b(w_pp_03_14), .i_c(w_pp_04_13), .ow_sum(w_sum_14), .ow_carry(w_carry_14));
wire w_sum_15, w_carry_15;
math_adder_carry_save CSA_15(.i_a(w_pp_05_12), .i_b(w_pp_06_11), .i_c(w_pp_07_10), .ow_sum(w_sum_15), .ow_carry(w_carry_15));
wire w_sum_16, w_carry_16;
math_adder_carry_save CSA_16(.i_a(w_pp_08_09), .i_b(w_pp_09_08), .i_c(w_pp_10_07), .ow_sum(w_sum_16), .ow_carry(w_carry_16));
wire w_sum_17, w_carry_17;
math_adder_carry_save CSA_17(.i_a(w_pp_03_15), .i_b(w_pp_04_14), .i_c(w_pp_05_13), .ow_sum(w_sum_17), .ow_carry(w_carry_17));
wire w_sum_18, w_carry_18;
math_adder_carry_save CSA_18(.i_a(w_pp_06_12), .i_b(w_pp_07_11), .i_c(w_pp_08_10), .ow_sum(w_sum_18), .ow_carry(w_carry_18));
wire w_sum_19, w_carry_19;
math_adder_carry_save CSA_19(.i_a(w_pp_04_15), .i_b(w_pp_05_14), .i_c(w_pp_06_13), .ow_sum(w_sum_19), .ow_carry(w_carry_19));
// Stage: 1, Max Height: 8
wire w_sum_20, w_carry_20;
math_adder_half HA_20(.i_a(w_pp_00_08), .i_b(w_pp_01_07), .ow_sum(w_sum_20), .ow_carry(w_carry_20));
wire w_sum_21, w_carry_21;
math_adder_carry_save CSA_21(.i_a(w_pp_00_09), .i_b(w_pp_01_08), .i_c(w_pp_02_07), .ow_sum(w_sum_21), .ow_carry(w_carry_21));
wire w_sum_22, w_carry_22;
math_adder_half HA_22(.i_a(w_pp_03_06), .i_b(w_pp_04_05), .ow_sum(w_sum_22), .ow_carry(w_carry_22));
wire w_sum_23, w_carry_23;
math_adder_carry_save CSA_23(.i_a(w_pp_00_10), .i_b(w_pp_01_09), .i_c(w_pp_02_08), .ow_sum(w_sum_23), .ow_carry(w_carry_23));
wire w_sum_24, w_carry_24;
math_adder_carry_save CSA_24(.i_a(w_pp_03_07), .i_b(w_pp_04_06), .i_c(w_pp_05_05), .ow_sum(w_sum_24), .ow_carry(w_carry_24));
wire w_sum_25, w_carry_25;
math_adder_half HA_25(.i_a(w_pp_06_04), .i_b(w_pp_07_03), .ow_sum(w_sum_25), .ow_carry(w_carry_25));
wire w_sum_26, w_carry_26;
math_adder_carry_save CSA_26(.i_a(w_pp_00_11), .i_b(w_pp_01_10), .i_c(w_pp_02_09), .ow_sum(w_sum_26), .ow_carry(w_carry_26));
wire w_sum_27, w_carry_27;
math_adder_carry_save CSA_27(.i_a(w_pp_03_08), .i_b(w_pp_04_07), .i_c(w_pp_05_06), .ow_sum(w_sum_27), .ow_carry(w_carry_27));
wire w_sum_28, w_carry_28;
math_adder_carry_save CSA_28(.i_a(w_pp_06_05), .i_b(w_pp_07_04), .i_c(w_pp_08_03), .ow_sum(w_sum_28), .ow_carry(w_carry_28));
wire w_sum_29, w_carry_29;
math_adder_half HA_29(.i_a(w_pp_09_02), .i_b(w_pp_10_01), .ow_sum(w_sum_29), .ow_carry(w_carry_29));
wire w_sum_30, w_carry_30;
math_adder_carry_save CSA_30(.i_a(w_pp_02_10), .i_b(w_pp_03_09), .i_c(w_pp_04_08), .ow_sum(w_sum_30), .ow_carry(w_carry_30));
wire w_sum_31, w_carry_31;
math_adder_carry_save CSA_31(.i_a(w_pp_05_07), .i_b(w_pp_06_06), .i_c(w_pp_07_05), .ow_sum(w_sum_31), .ow_carry(w_carry_31));
wire w_sum_32, w_carry_32;
math_adder_carry_save CSA_32(.i_a(w_pp_08_04), .i_b(w_pp_09_03), .i_c(w_pp_10_02), .ow_sum(w_sum_32), .ow_carry(w_carry_32));
wire w_sum_33, w_carry_33;
math_adder_carry_save CSA_33(.i_a(w_pp_11_01), .i_b(w_pp_12_00), .i_c(w_sum_0), .ow_sum(w_sum_33), .ow_carry(w_carry_33));
wire w_sum_34, w_carry_34;
math_adder_carry_save CSA_34(.i_a(w_pp_05_08), .i_b(w_pp_06_07), .i_c(w_pp_07_06), .ow_sum(w_sum_34), .ow_carry(w_carry_34));
wire w_sum_35, w_carry_35;
math_adder_carry_save CSA_35(.i_a(w_pp_08_05), .i_b(w_pp_09_04), .i_c(w_pp_10_03), .ow_sum(w_sum_35), .ow_carry(w_carry_35));
wire w_sum_36, w_carry_36;
math_adder_carry_save CSA_36(.i_a(w_pp_11_02), .i_b(w_pp_12_01), .i_c(w_pp_13_00), .ow_sum(w_sum_36), .ow_carry(w_carry_36));
wire w_sum_37, w_carry_37;
math_adder_carry_save CSA_37(.i_a(w_carry_0), .i_b(w_sum_1), .i_c(w_sum_2), .ow_sum(w_sum_37), .ow_carry(w_carry_37));
wire w_sum_38, w_carry_38;
math_adder_carry_save CSA_38(.i_a(w_pp_08_06), .i_b(w_pp_09_05), .i_c(w_pp_10_04), .ow_sum(w_sum_38), .ow_carry(w_carry_38));
wire w_sum_39, w_carry_39;
math_adder_carry_save CSA_39(.i_a(w_pp_11_03), .i_b(w_pp_12_02), .i_c(w_pp_13_01), .ow_sum(w_sum_39), .ow_carry(w_carry_39));
wire w_sum_40, w_carry_40;
math_adder_carry_save CSA_40(.i_a(w_pp_14_00), .i_b(w_carry_1), .i_c(w_carry_2), .ow_sum(w_sum_40), .ow_carry(w_carry_40));
wire w_sum_41, w_carry_41;
math_adder_carry_save CSA_41(.i_a(w_sum_3), .i_b(w_sum_4), .i_c(w_sum_5), .ow_sum(w_sum_41), .ow_carry(w_carry_41));
wire w_sum_42, w_carry_42;
math_adder_carry_save CSA_42(.i_a(w_pp_11_04), .i_b(w_pp_12_03), .i_c(w_pp_13_02), .ow_sum(w_sum_42), .ow_carry(w_carry_42));
wire w_sum_43, w_carry_43;
math_adder_carry_save CSA_43(.i_a(w_pp_14_01), .i_b(w_pp_15_00), .i_c(w_carry_3), .ow_sum(w_sum_43), .ow_carry(w_carry_43));
wire w_sum_44, w_carry_44;
math_adder_carry_save CSA_44(.i_a(w_carry_4), .i_b(w_carry_5), .i_c(w_sum_6), .ow_sum(w_sum_44), .ow_carry(w_carry_44));
wire w_sum_45, w_carry_45;
math_adder_carry_save CSA_45(.i_a(w_sum_7), .i_b(w_sum_8), .i_c(w_sum_9), .ow_sum(w_sum_45), .ow_carry(w_carry_45));
wire w_sum_46, w_carry_46;
math_adder_carry_save CSA_46(.i_a(w_pp_12_04), .i_b(w_pp_13_03), .i_c(w_pp_14_02), .ow_sum(w_sum_46), .ow_carry(w_carry_46));
wire w_sum_47, w_carry_47;
math_adder_carry_save CSA_47(.i_a(w_pp_15_01), .i_b(w_carry_6), .i_c(w_carry_7), .ow_sum(w_sum_47), .ow_carry(w_carry_47));
wire w_sum_48, w_carry_48;
math_adder_carry_save CSA_48(.i_a(w_carry_8), .i_b(w_carry_9), .i_c(w_sum_10), .ow_sum(w_sum_48), .ow_carry(w_carry_48));
wire w_sum_49, w_carry_49;
math_adder_carry_save CSA_49(.i_a(w_sum_11), .i_b(w_sum_12), .i_c(w_sum_13), .ow_sum(w_sum_49), .ow_carry(w_carry_49));
wire w_sum_50, w_carry_50;
math_adder_carry_save CSA_50(.i_a(w_pp_11_06), .i_b(w_pp_12_05), .i_c(w_pp_13_04), .ow_sum(w_sum_50), .ow_carry(w_carry_50));
wire w_sum_51, w_carry_51;
math_adder_carry_save CSA_51(.i_a(w_pp_14_03), .i_b(w_pp_15_02), .i_c(w_carry_10), .ow_sum(w_sum_51), .ow_carry(w_carry_51));
wire w_sum_52, w_carry_52;
math_adder_carry_save CSA_52(.i_a(w_carry_11), .i_b(w_carry_12), .i_c(w_carry_13), .ow_sum(w_sum_52), .ow_carry(w_carry_52));
wire w_sum_53, w_carry_53;
math_adder_carry_save CSA_53(.i_a(w_sum_14), .i_b(w_sum_15), .i_c(w_sum_16), .ow_sum(w_sum_53), .ow_carry(w_carry_53));
wire w_sum_54, w_carry_54;
math_adder_carry_save CSA_54(.i_a(w_pp_09_09), .i_b(w_pp_10_08), .i_c(w_pp_11_07), .ow_sum(w_sum_54), .ow_carry(w_carry_54));
wire w_sum_55, w_carry_55;
math_adder_carry_save CSA_55(.i_a(w_pp_12_06), .i_b(w_pp_13_05), .i_c(w_pp_14_04), .ow_sum(w_sum_55), .ow_carry(w_carry_55));
wire w_sum_56, w_carry_56;
math_adder_carry_save CSA_56(.i_a(w_pp_15_03), .i_b(w_carry_14), .i_c(w_carry_15), .ow_sum(w_sum_56), .ow_carry(w_carry_56));
wire w_sum_57, w_carry_57;
math_adder_carry_save CSA_57(.i_a(w_carry_16), .i_b(w_sum_17), .i_c(w_sum_18), .ow_sum(w_sum_57), .ow_carry(w_carry_57));
wire w_sum_58, w_carry_58;
math_adder_carry_save CSA_58(.i_a(w_pp_07_12), .i_b(w_pp_08_11), .i_c(w_pp_09_10), .ow_sum(w_sum_58), .ow_carry(w_carry_58));
wire w_sum_59, w_carry_59;
math_adder_carry_save CSA_59(.i_a(w_pp_10_09), .i_b(w_pp_11_08), .i_c(w_pp_12_07), .ow_sum(w_sum_59), .ow_carry(w_carry_59));
wire w_sum_60, w_carry_60;
math_adder_carry_save CSA_60(.i_a(w_pp_13_06), .i_b(w_pp_14_05), .i_c(w_pp_15_04), .ow_sum(w_sum_60), .ow_carry(w_carry_60));
wire w_sum_61, w_carry_61;
math_adder_carry_save CSA_61(.i_a(w_carry_17), .i_b(w_carry_18), .i_c(w_sum_19), .ow_sum(w_sum_61), .ow_carry(w_carry_61));
wire w_sum_62, w_carry_62;
math_adder_carry_save CSA_62(.i_a(w_pp_05_15), .i_b(w_pp_06_14), .i_c(w_pp_07_13), .ow_sum(w_sum_62), .ow_carry(w_carry_62));
wire w_sum_63, w_carry_63;
math_adder_carry_save CSA_63(.i_a(w_pp_08_12), .i_b(w_pp_09_11), .i_c(w_pp_10_10), .ow_sum(w_sum_63), .ow_carry(w_carry_63));
wire w_sum_64, w_carry_64;
math_adder_carry_save CSA_64(.i_a(w_pp_11_09), .i_b(w_pp_12_08), .i_c(w_pp_13_07), .ow_sum(w_sum_64), .ow_carry(w_carry_64));
wire w_sum_65, w_carry_65;
math_adder_carry_save CSA_65(.i_a(w_pp_14_06), .i_b(w_pp_15_05), .i_c(w_carry_19), .ow_sum(w_sum_65), .ow_carry(w_carry_65));
wire w_sum_66, w_carry_66;
math_adder_carry_save CSA_66(.i_a(w_pp_06_15), .i_b(w_pp_07_14), .i_c(w_pp_08_13), .ow_sum(w_sum_66), .ow_carry(w_carry_66));
wire w_sum_67, w_carry_67;
math_adder_carry_save CSA_67(.i_a(w_pp_09_12), .i_b(w_pp_10_11), .i_c(w_pp_11_10), .ow_sum(w_sum_67), .ow_carry(w_carry_67));
wire w_sum_68, w_carry_68;
math_adder_carry_save CSA_68(.i_a(w_pp_12_09), .i_b(w_pp_13_08), .i_c(w_pp_14_07), .ow_sum(w_sum_68), .ow_carry(w_carry_68));
wire w_sum_69, w_carry_69;
math_adder_carry_save CSA_69(.i_a(w_pp_07_15), .i_b(w_pp_08_14), .i_c(w_pp_09_13), .ow_sum(w_sum_69), .ow_carry(w_carry_69));
wire w_sum_70, w_carry_70;
math_adder_carry_save CSA_70(.i_a(w_pp_10_12), .i_b(w_pp_11_11), .i_c(w_pp_12_10), .ow_sum(w_sum_70), .ow_carry(w_carry_70));
wire w_sum_71, w_carry_71;
math_adder_carry_save CSA_71(.i_a(w_pp_08_15), .i_b(w_pp_09_14), .i_c(w_pp_10_13), .ow_sum(w_sum_71), .ow_carry(w_carry_71));
// Stage: 2, Max Height: 6
wire w_sum_72, w_carry_72;
math_adder_half HA_72(.i_a(w_pp_00_06), .i_b(w_pp_01_05), .ow_sum(w_sum_72), .ow_carry(w_carry_72));
wire w_sum_73, w_carry_73;
math_adder_carry_save CSA_73(.i_a(w_pp_00_07), .i_b(w_pp_01_06), .i_c(w_pp_02_05), .ow_sum(w_sum_73), .ow_carry(w_carry_73));
wire w_sum_74, w_carry_74;
math_adder_half HA_74(.i_a(w_pp_03_04), .i_b(w_pp_04_03), .ow_sum(w_sum_74), .ow_carry(w_carry_74));
wire w_sum_75, w_carry_75;
math_adder_carry_save CSA_75(.i_a(w_pp_02_06), .i_b(w_pp_03_05), .i_c(w_pp_04_04), .ow_sum(w_sum_75), .ow_carry(w_carry_75));
wire w_sum_76, w_carry_76;
math_adder_carry_save CSA_76(.i_a(w_pp_05_03), .i_b(w_pp_06_02), .i_c(w_pp_07_01), .ow_sum(w_sum_76), .ow_carry(w_carry_76));
wire w_sum_77, w_carry_77;
math_adder_carry_save CSA_77(.i_a(w_pp_05_04), .i_b(w_pp_06_03), .i_c(w_pp_07_02), .ow_sum(w_sum_77), .ow_carry(w_carry_77));
wire w_sum_78, w_carry_78;
math_adder_carry_save CSA_78(.i_a(w_pp_08_01), .i_b(w_pp_09_00), .i_c(w_carry_20), .ow_sum(w_sum_78), .ow_carry(w_carry_78));
wire w_sum_79, w_carry_79;
math_adder_carry_save CSA_79(.i_a(w_pp_08_02), .i_b(w_pp_09_01), .i_c(w_pp_10_00), .ow_sum(w_sum_79), .ow_carry(w_carry_79));
wire w_sum_80, w_carry_80;
math_adder_carry_save CSA_80(.i_a(w_carry_21), .i_b(w_carry_22), .i_c(w_sum_23), .ow_sum(w_sum_80), .ow_carry(w_carry_80));
wire w_sum_81, w_carry_81;
math_adder_carry_save CSA_81(.i_a(w_pp_11_00), .i_b(w_carry_23), .i_c(w_carry_24), .ow_sum(w_sum_81), .ow_carry(w_carry_81));
wire w_sum_82, w_carry_82;
math_adder_carry_save CSA_82(.i_a(w_carry_25), .i_b(w_sum_26), .i_c(w_sum_27), .ow_sum(w_sum_82), .ow_carry(w_carry_82));
wire w_sum_83, w_carry_83;
math_adder_carry_save CSA_83(.i_a(w_carry_26), .i_b(w_carry_27), .i_c(w_carry_28), .ow_sum(w_sum_83), .ow_carry(w_carry_83));
wire w_sum_84, w_carry_84;
math_adder_carry_save CSA_84(.i_a(w_carry_29), .i_b(w_sum_30), .i_c(w_sum_31), .ow_sum(w_sum_84), .ow_carry(w_carry_84));
wire w_sum_85, w_carry_85;
math_adder_carry_save CSA_85(.i_a(w_carry_30), .i_b(w_carry_31), .i_c(w_carry_32), .ow_sum(w_sum_85), .ow_carry(w_carry_85));
wire w_sum_86, w_carry_86;
math_adder_carry_save CSA_86(.i_a(w_carry_33), .i_b(w_sum_34), .i_c(w_sum_35), .ow_sum(w_sum_86), .ow_carry(w_carry_86));
wire w_sum_87, w_carry_87;
math_adder_carry_save CSA_87(.i_a(w_carry_34), .i_b(w_carry_35), .i_c(w_carry_36), .ow_sum(w_sum_87), .ow_carry(w_carry_87));
wire w_sum_88, w_carry_88;
math_adder_carry_save CSA_88(.i_a(w_carry_37), .i_b(w_sum_38), .i_c(w_sum_39), .ow_sum(w_sum_88), .ow_carry(w_carry_88));
wire w_sum_89, w_carry_89;
math_adder_carry_save CSA_89(.i_a(w_carry_38), .i_b(w_carry_39), .i_c(w_carry_40), .ow_sum(w_sum_89), .ow_carry(w_carry_89));
wire w_sum_90, w_carry_90;
math_adder_carry_save CSA_90(.i_a(w_carry_41), .i_b(w_sum_42), .i_c(w_sum_43), .ow_sum(w_sum_90), .ow_carry(w_carry_90));
wire w_sum_91, w_carry_91;
math_adder_carry_save CSA_91(.i_a(w_carry_42), .i_b(w_carry_43), .i_c(w_carry_44), .ow_sum(w_sum_91), .ow_carry(w_carry_91));
wire w_sum_92, w_carry_92;
math_adder_carry_save CSA_92(.i_a(w_carry_45), .i_b(w_sum_46), .i_c(w_sum_47), .ow_sum(w_sum_92), .ow_carry(w_carry_92));
wire w_sum_93, w_carry_93;
math_adder_carry_save CSA_93(.i_a(w_carry_46), .i_b(w_carry_47), .i_c(w_carry_48), .ow_sum(w_sum_93), .ow_carry(w_carry_93));
wire w_sum_94, w_carry_94;
math_adder_carry_save CSA_94(.i_a(w_carry_49), .i_b(w_sum_50), .i_c(w_sum_51), .ow_sum(w_sum_94), .ow_carry(w_carry_94));
wire w_sum_95, w_carry_95;
math_adder_carry_save CSA_95(.i_a(w_carry_50), .i_b(w_carry_51), .i_c(w_carry_52), .ow_sum(w_sum_95), .ow_carry(w_carry_95));
wire w_sum_96, w_carry_96;
math_adder_carry_save CSA_96(.i_a(w_carry_53), .i_b(w_sum_54), .i_c(w_sum_55), .ow_sum(w_sum_96), .ow_carry(w_carry_96));
wire w_sum_97, w_carry_97;
math_adder_carry_save CSA_97(.i_a(w_carry_54), .i_b(w_carry_55), .i_c(w_carry_56), .ow_sum(w_sum_97), .ow_carry(w_carry_97));
wire w_sum_98, w_carry_98;
math_adder_carry_save CSA_98(.i_a(w_carry_57), .i_b(w_sum_58), .i_c(w_sum_59), .ow_sum(w_sum_98), .ow_carry(w_carry_98));
wire w_sum_99, w_carry_99;
math_adder_carry_save CSA_99(.i_a(w_carry_58), .i_b(w_carry_59), .i_c(w_carry_60), .ow_sum(w_sum_99), .ow_carry(w_carry_99));
wire w_sum_100, w_carry_100;
math_adder_carry_save CSA_100(.i_a(w_carry_61), .i_b(w_sum_62), .i_c(w_sum_63), .ow_sum(w_sum_100), .ow_carry(w_carry_100));
wire w_sum_101, w_carry_101;
math_adder_carry_save CSA_101(.i_a(w_pp_15_06), .i_b(w_carry_62), .i_c(w_carry_63), .ow_sum(w_sum_101), .ow_carry(w_carry_101));
wire w_sum_102, w_carry_102;
math_adder_carry_save CSA_102(.i_a(w_carry_64), .i_b(w_carry_65), .i_c(w_sum_66), .ow_sum(w_sum_102), .ow_carry(w_carry_102));
wire w_sum_103, w_carry_103;
math_adder_carry_save CSA_103(.i_a(w_pp_13_09), .i_b(w_pp_14_08), .i_c(w_pp_15_07), .ow_sum(w_sum_103), .ow_carry(w_carry_103));
wire w_sum_104, w_carry_104;
math_adder_carry_save CSA_104(.i_a(w_carry_66), .i_b(w_carry_67), .i_c(w_carry_68), .ow_sum(w_sum_104), .ow_carry(w_carry_104));
wire w_sum_105, w_carry_105;
math_adder_carry_save CSA_105(.i_a(w_pp_11_12), .i_b(w_pp_12_11), .i_c(w_pp_13_10), .ow_sum(w_sum_105), .ow_carry(w_carry_105));
wire w_sum_106, w_carry_106;
math_adder_carry_save CSA_106(.i_a(w_pp_14_09), .i_b(w_pp_15_08), .i_c(w_carry_69), .ow_sum(w_sum_106), .ow_carry(w_carry_106));
wire w_sum_107, w_carry_107;
math_adder_carry_save CSA_107(.i_a(w_pp_09_15), .i_b(w_pp_10_14), .i_c(w_pp_11_13), .ow_sum(w_sum_107), .ow_carry(w_carry_107));
wire w_sum_108, w_carry_108;
math_adder_carry_save CSA_108(.i_a(w_pp_12_12), .i_b(w_pp_13_11), .i_c(w_pp_14_10), .ow_sum(w_sum_108), .ow_carry(w_carry_108));
wire w_sum_109, w_carry_109;
math_adder_carry_save CSA_109(.i_a(w_pp_10_15), .i_b(w_pp_11_14), .i_c(w_pp_12_13), .ow_sum(w_sum_109), .ow_carry(w_carry_109));
// Stage: 3, Max Height: 4
wire w_sum_110, w_carry_110;
math_adder_half HA_110(.i_a(w_pp_00_04), .i_b(w_pp_01_03), .ow_sum(w_sum_110), .ow_carry(w_carry_110));
wire w_sum_111, w_carry_111;
math_adder_carry_save CSA_111(.i_a(w_pp_00_05), .i_b(w_pp_01_04), .i_c(w_pp_02_03), .ow_sum(w_sum_111), .ow_carry(w_carry_111));
wire w_sum_112, w_carry_112;
math_adder_half HA_112(.i_a(w_pp_03_02), .i_b(w_pp_04_01), .ow_sum(w_sum_112), .ow_carry(w_carry_112));
wire w_sum_113, w_carry_113;
math_adder_carry_save CSA_113(.i_a(w_pp_02_04), .i_b(w_pp_03_03), .i_c(w_pp_04_02), .ow_sum(w_sum_113), .ow_carry(w_carry_113));
wire w_sum_114, w_carry_114;
math_adder_carry_save CSA_114(.i_a(w_pp_05_01), .i_b(w_pp_06_00), .i_c(w_sum_72), .ow_sum(w_sum_114), .ow_carry(w_carry_114));
wire w_sum_115, w_carry_115;
math_adder_carry_save CSA_115(.i_a(w_pp_05_02), .i_b(w_pp_06_01), .i_c(w_pp_07_00), .ow_sum(w_sum_115), .ow_carry(w_carry_115));
wire w_sum_116, w_carry_116;
math_adder_carry_save CSA_116(.i_a(w_carry_72), .i_b(w_sum_73), .i_c(w_sum_74), .ow_sum(w_sum_116), .ow_carry(w_carry_116));
wire w_sum_117, w_carry_117;
math_adder_carry_save CSA_117(.i_a(w_pp_08_00), .i_b(w_sum_20), .i_c(w_carry_73), .ow_sum(w_sum_117), .ow_carry(w_carry_117));
wire w_sum_118, w_carry_118;
math_adder_carry_save CSA_118(.i_a(w_carry_74), .i_b(w_sum_75), .i_c(w_sum_76), .ow_sum(w_sum_118), .ow_carry(w_carry_118));
wire w_sum_119, w_carry_119;
math_adder_carry_save CSA_119(.i_a(w_sum_21), .i_b(w_sum_22), .i_c(w_carry_75), .ow_sum(w_sum_119), .ow_carry(w_carry_119));
wire w_sum_120, w_carry_120;
math_adder_carry_save CSA_120(.i_a(w_carry_76), .i_b(w_sum_77), .i_c(w_sum_78), .ow_sum(w_sum_120), .ow_carry(w_carry_120));
wire w_sum_121, w_carry_121;
math_adder_carry_save CSA_121(.i_a(w_sum_24), .i_b(w_sum_25), .i_c(w_carry_77), .ow_sum(w_sum_121), .ow_carry(w_carry_121));
wire w_sum_122, w_carry_122;
math_adder_carry_save CSA_122(.i_a(w_carry_78), .i_b(w_sum_79), .i_c(w_sum_80), .ow_sum(w_sum_122), .ow_carry(w_carry_122));
wire w_sum_123, w_carry_123;
math_adder_carry_save CSA_123(.i_a(w_sum_28), .i_b(w_sum_29), .i_c(w_carry_79), .ow_sum(w_sum_123), .ow_carry(w_carry_123));
wire w_sum_124, w_carry_124;
math_adder_carry_save CSA_124(.i_a(w_carry_80), .i_b(w_sum_81), .i_c(w_sum_82), .ow_sum(w_sum_124), .ow_carry(w_carry_124));
wire w_sum_125, w_carry_125;
math_adder_carry_save CSA_125(.i_a(w_sum_32), .i_b(w_sum_33), .i_c(w_carry_81), .ow_sum(w_sum_125), .ow_carry(w_carry_125));
wire w_sum_126, w_carry_126;
math_adder_carry_save CSA_126(.i_a(w_carry_82), .i_b(w_sum_83), .i_c(w_sum_84), .ow_sum(w_sum_126), .ow_carry(w_carry_126));
wire w_sum_127, w_carry_127;
math_adder_carry_save CSA_127(.i_a(w_sum_36), .i_b(w_sum_37), .i_c(w_carry_83), .ow_sum(w_sum_127), .ow_carry(w_carry_127));
wire w_sum_128, w_carry_128;
math_adder_carry_save CSA_128(.i_a(w_carry_84), .i_b(w_sum_85), .i_c(w_sum_86), .ow_sum(w_sum_128), .ow_carry(w_carry_128));
wire w_sum_129, w_carry_129;
math_adder_carry_save CSA_129(.i_a(w_sum_40), .i_b(w_sum_41), .i_c(w_carry_85), .ow_sum(w_sum_129), .ow_carry(w_carry_129));
wire w_sum_130, w_carry_130;
math_adder_carry_save CSA_130(.i_a(w_carry_86), .i_b(w_sum_87), .i_c(w_sum_88), .ow_sum(w_sum_130), .ow_carry(w_carry_130));
wire w_sum_131, w_carry_131;
math_adder_carry_save CSA_131(.i_a(w_sum_44), .i_b(w_sum_45), .i_c(w_carry_87), .ow_sum(w_sum_131), .ow_carry(w_carry_131));
wire w_sum_132, w_carry_132;
math_adder_carry_save CSA_132(.i_a(w_carry_88), .i_b(w_sum_89), .i_c(w_sum_90), .ow_sum(w_sum_132), .ow_carry(w_carry_132));
wire w_sum_133, w_carry_133;
math_adder_carry_save CSA_133(.i_a(w_sum_48), .i_b(w_sum_49), .i_c(w_carry_89), .ow_sum(w_sum_133), .ow_carry(w_carry_133));
wire w_sum_134, w_carry_134;
math_adder_carry_save CSA_134(.i_a(w_carry_90), .i_b(w_sum_91), .i_c(w_sum_92), .ow_sum(w_sum_134), .ow_carry(w_carry_134));
wire w_sum_135, w_carry_135;
math_adder_carry_save CSA_135(.i_a(w_sum_52), .i_b(w_sum_53), .i_c(w_carry_91), .ow_sum(w_sum_135), .ow_carry(w_carry_135));
wire w_sum_136, w_carry_136;
math_adder_carry_save CSA_136(.i_a(w_carry_92), .i_b(w_sum_93), .i_c(w_sum_94), .ow_sum(w_sum_136), .ow_carry(w_carry_136));
wire w_sum_137, w_carry_137;
math_adder_carry_save CSA_137(.i_a(w_sum_56), .i_b(w_sum_57), .i_c(w_carry_93), .ow_sum(w_sum_137), .ow_carry(w_carry_137));
wire w_sum_138, w_carry_138;
math_adder_carry_save CSA_138(.i_a(w_carry_94), .i_b(w_sum_95), .i_c(w_sum_96), .ow_sum(w_sum_138), .ow_carry(w_carry_138));
wire w_sum_139, w_carry_139;
math_adder_carry_save CSA_139(.i_a(w_sum_60), .i_b(w_sum_61), .i_c(w_carry_95), .ow_sum(w_sum_139), .ow_carry(w_carry_139));
wire w_sum_140, w_carry_140;
math_adder_carry_save CSA_140(.i_a(w_carry_96), .i_b(w_sum_97), .i_c(w_sum_98), .ow_sum(w_sum_140), .ow_carry(w_carry_140));
wire w_sum_141, w_carry_141;
math_adder_carry_save CSA_141(.i_a(w_sum_64), .i_b(w_sum_65), .i_c(w_carry_97), .ow_sum(w_sum_141), .ow_carry(w_carry_141));
wire w_sum_142, w_carry_142;
math_adder_carry_save CSA_142(.i_a(w_carry_98), .i_b(w_sum_99), .i_c(w_sum_100), .ow_sum(w_sum_142), .ow_carry(w_carry_142));
wire w_sum_143, w_carry_143;
math_adder_carry_save CSA_143(.i_a(w_sum_67), .i_b(w_sum_68), .i_c(w_carry_99), .ow_sum(w_sum_143), .ow_carry(w_carry_143));
wire w_sum_144, w_carry_144;
math_adder_carry_save CSA_144(.i_a(w_carry_100), .i_b(w_sum_101), .i_c(w_sum_102), .ow_sum(w_sum_144), .ow_carry(w_carry_144));
wire w_sum_145, w_carry_145;
math_adder_carry_save CSA_145(.i_a(w_sum_69), .i_b(w_sum_70), .i_c(w_carry_101), .ow_sum(w_sum_145), .ow_carry(w_carry_145));
wire w_sum_146, w_carry_146;
math_adder_carry_save CSA_146(.i_a(w_carry_102), .i_b(w_sum_103), .i_c(w_sum_104), .ow_sum(w_sum_146), .ow_carry(w_carry_146));
wire w_sum_147, w_carry_147;
math_adder_carry_save CSA_147(.i_a(w_carry_70), .i_b(w_sum_71), .i_c(w_carry_103), .ow_sum(w_sum_147), .ow_carry(w_carry_147));
wire w_sum_148, w_carry_148;
math_adder_carry_save CSA_148(.i_a(w_carry_104), .i_b(w_sum_105), .i_c(w_sum_106), .ow_sum(w_sum_148), .ow_carry(w_carry_148));
wire w_sum_149, w_carry_149;
math_adder_carry_save CSA_149(.i_a(w_pp_15_09), .i_b(w_carry_71), .i_c(w_carry_105), .ow_sum(w_sum_149), .ow_carry(w_carry_149));
wire w_sum_150, w_carry_150;
math_adder_carry_save CSA_150(.i_a(w_carry_106), .i_b(w_sum_107), .i_c(w_sum_108), .ow_sum(w_sum_150), .ow_carry(w_carry_150));
wire w_sum_151, w_carry_151;
math_adder_carry_save CSA_151(.i_a(w_pp_13_12), .i_b(w_pp_14_11), .i_c(w_pp_15_10), .ow_sum(w_sum_151), .ow_carry(w_carry_151));
wire w_sum_152, w_carry_152;
math_adder_carry_save CSA_152(.i_a(w_carry_107), .i_b(w_carry_108), .i_c(w_sum_109), .ow_sum(w_sum_152), .ow_carry(w_carry_152));
wire w_sum_153, w_carry_153;
math_adder_carry_save CSA_153(.i_a(w_pp_11_15), .i_b(w_pp_12_14), .i_c(w_pp_13_13), .ow_sum(w_sum_153), .ow_carry(w_carry_153));
wire w_sum_154, w_carry_154;
math_adder_carry_save CSA_154(.i_a(w_pp_14_12), .i_b(w_pp_15_11), .i_c(w_carry_109), .ow_sum(w_sum_154), .ow_carry(w_carry_154));
wire w_sum_155, w_carry_155;
math_adder_carry_save CSA_155(.i_a(w_pp_12_15), .i_b(w_pp_13_14), .i_c(w_pp_14_13), .ow_sum(w_sum_155), .ow_carry(w_carry_155));
// Stage: 4, Max Height: 3
wire w_sum_156, w_carry_156;
math_adder_half HA_156(.i_a(w_pp_00_03), .i_b(w_pp_01_02), .ow_sum(w_sum_156), .ow_carry(w_carry_156));
wire w_sum_157, w_carry_157;
math_adder_carry_save CSA_157(.i_a(w_pp_02_02), .i_b(w_pp_03_01), .i_c(w_pp_04_00), .ow_sum(w_sum_157), .ow_carry(w_carry_157));
wire w_sum_158, w_carry_158;
math_adder_carry_save CSA_158(.i_a(w_pp_05_00), .i_b(w_carry_110), .i_c(w_sum_111), .ow_sum(w_sum_158), .ow_carry(w_carry_158));
wire w_sum_159, w_carry_159;
math_adder_carry_save CSA_159(.i_a(w_carry_111), .i_b(w_carry_112), .i_c(w_sum_113), .ow_sum(w_sum_159), .ow_carry(w_carry_159));
wire w_sum_160, w_carry_160;
math_adder_carry_save CSA_160(.i_a(w_carry_113), .i_b(w_carry_114), .i_c(w_sum_115), .ow_sum(w_sum_160), .ow_carry(w_carry_160));
wire w_sum_161, w_carry_161;
math_adder_carry_save CSA_161(.i_a(w_carry_115), .i_b(w_carry_116), .i_c(w_sum_117), .ow_sum(w_sum_161), .ow_carry(w_carry_161));
wire w_sum_162, w_carry_162;
math_adder_carry_save CSA_162(.i_a(w_carry_117), .i_b(w_carry_118), .i_c(w_sum_119), .ow_sum(w_sum_162), .ow_carry(w_carry_162));
wire w_sum_163, w_carry_163;
math_adder_carry_save CSA_163(.i_a(w_carry_119), .i_b(w_carry_120), .i_c(w_sum_121), .ow_sum(w_sum_163), .ow_carry(w_carry_163));
wire w_sum_164, w_carry_164;
math_adder_carry_save CSA_164(.i_a(w_carry_121), .i_b(w_carry_122), .i_c(w_sum_123), .ow_sum(w_sum_164), .ow_carry(w_carry_164));
wire w_sum_165, w_carry_165;
math_adder_carry_save CSA_165(.i_a(w_carry_123), .i_b(w_carry_124), .i_c(w_sum_125), .ow_sum(w_sum_165), .ow_carry(w_carry_165));
wire w_sum_166, w_carry_166;
math_adder_carry_save CSA_166(.i_a(w_carry_125), .i_b(w_carry_126), .i_c(w_sum_127), .ow_sum(w_sum_166), .ow_carry(w_carry_166));
wire w_sum_167, w_carry_167;
math_adder_carry_save CSA_167(.i_a(w_carry_127), .i_b(w_carry_128), .i_c(w_sum_129), .ow_sum(w_sum_167), .ow_carry(w_carry_167));
wire w_sum_168, w_carry_168;
math_adder_carry_save CSA_168(.i_a(w_carry_129), .i_b(w_carry_130), .i_c(w_sum_131), .ow_sum(w_sum_168), .ow_carry(w_carry_168));
wire w_sum_169, w_carry_169;
math_adder_carry_save CSA_169(.i_a(w_carry_131), .i_b(w_carry_132), .i_c(w_sum_133), .ow_sum(w_sum_169), .ow_carry(w_carry_169));
wire w_sum_170, w_carry_170;
math_adder_carry_save CSA_170(.i_a(w_carry_133), .i_b(w_carry_134), .i_c(w_sum_135), .ow_sum(w_sum_170), .ow_carry(w_carry_170));
wire w_sum_171, w_carry_171;
math_adder_carry_save CSA_171(.i_a(w_carry_135), .i_b(w_carry_136), .i_c(w_sum_137), .ow_sum(w_sum_171), .ow_carry(w_carry_171));
wire w_sum_172, w_carry_172;
math_adder_carry_save CSA_172(.i_a(w_carry_137), .i_b(w_carry_138), .i_c(w_sum_139), .ow_sum(w_sum_172), .ow_carry(w_carry_172));
wire w_sum_173, w_carry_173;
math_adder_carry_save CSA_173(.i_a(w_carry_139), .i_b(w_carry_140), .i_c(w_sum_141), .ow_sum(w_sum_173), .ow_carry(w_carry_173));
wire w_sum_174, w_carry_174;
math_adder_carry_save CSA_174(.i_a(w_carry_141), .i_b(w_carry_142), .i_c(w_sum_143), .ow_sum(w_sum_174), .ow_carry(w_carry_174));
wire w_sum_175, w_carry_175;
math_adder_carry_save CSA_175(.i_a(w_carry_143), .i_b(w_carry_144), .i_c(w_sum_145), .ow_sum(w_sum_175), .ow_carry(w_carry_175));
wire w_sum_176, w_carry_176;
math_adder_carry_save CSA_176(.i_a(w_carry_145), .i_b(w_carry_146), .i_c(w_sum_147), .ow_sum(w_sum_176), .ow_carry(w_carry_176));
wire w_sum_177, w_carry_177;
math_adder_carry_save CSA_177(.i_a(w_carry_147), .i_b(w_carry_148), .i_c(w_sum_149), .ow_sum(w_sum_177), .ow_carry(w_carry_177));
wire w_sum_178, w_carry_178;
math_adder_carry_save CSA_178(.i_a(w_carry_149), .i_b(w_carry_150), .i_c(w_sum_151), .ow_sum(w_sum_178), .ow_carry(w_carry_178));
wire w_sum_179, w_carry_179;
math_adder_carry_save CSA_179(.i_a(w_carry_151), .i_b(w_carry_152), .i_c(w_sum_153), .ow_sum(w_sum_179), .ow_carry(w_carry_179));
wire w_sum_180, w_carry_180;
math_adder_carry_save CSA_180(.i_a(w_pp_15_12), .i_b(w_carry_153), .i_c(w_carry_154), .ow_sum(w_sum_180), .ow_carry(w_carry_180));
wire w_sum_181, w_carry_181;
math_adder_carry_save CSA_181(.i_a(w_pp_13_15), .i_b(w_pp_14_14), .i_c(w_pp_15_13), .ow_sum(w_sum_181), .ow_carry(w_carry_181));
// Stage: 5, Max Height: 2
wire w_sum_182, w_carry_182;
math_adder_half HA_182(.i_a(w_pp_00_02), .i_b(w_pp_01_01), .ow_sum(w_sum_182), .ow_carry(w_carry_182));
wire w_sum_183, w_carry_183;
math_adder_carry_save CSA_183(.i_a(w_pp_02_01), .i_b(w_pp_03_00), .i_c(w_sum_156), .ow_sum(w_sum_183), .ow_carry(w_carry_183));
wire w_sum_184, w_carry_184;
math_adder_carry_save CSA_184(.i_a(w_sum_110), .i_b(w_carry_156), .i_c(w_sum_157), .ow_sum(w_sum_184), .ow_carry(w_carry_184));
wire w_sum_185, w_carry_185;
math_adder_carry_save CSA_185(.i_a(w_sum_112), .i_b(w_carry_157), .i_c(w_sum_158), .ow_sum(w_sum_185), .ow_carry(w_carry_185));
wire w_sum_186, w_carry_186;
math_adder_carry_save CSA_186(.i_a(w_sum_114), .i_b(w_carry_158), .i_c(w_sum_159), .ow_sum(w_sum_186), .ow_carry(w_carry_186));
wire w_sum_187, w_carry_187;
math_adder_carry_save CSA_187(.i_a(w_sum_116), .i_b(w_carry_159), .i_c(w_sum_160), .ow_sum(w_sum_187), .ow_carry(w_carry_187));
wire w_sum_188, w_carry_188;
math_adder_carry_save CSA_188(.i_a(w_sum_118), .i_b(w_carry_160), .i_c(w_sum_161), .ow_sum(w_sum_188), .ow_carry(w_carry_188));
wire w_sum_189, w_carry_189;
math_adder_carry_save CSA_189(.i_a(w_sum_120), .i_b(w_carry_161), .i_c(w_sum_162), .ow_sum(w_sum_189), .ow_carry(w_carry_189));
wire w_sum_190, w_carry_190;
math_adder_carry_save CSA_190(.i_a(w_sum_122), .i_b(w_carry_162), .i_c(w_sum_163), .ow_sum(w_sum_190), .ow_carry(w_carry_190));
wire w_sum_191, w_carry_191;
math_adder_carry_save CSA_191(.i_a(w_sum_124), .i_b(w_carry_163), .i_c(w_sum_164), .ow_sum(w_sum_191), .ow_carry(w_carry_191));
wire w_sum_192, w_carry_192;
math_adder_carry_save CSA_192(.i_a(w_sum_126), .i_b(w_carry_164), .i_c(w_sum_165), .ow_sum(w_sum_192), .ow_carry(w_carry_192));
wire w_sum_193, w_carry_193;
math_adder_carry_save CSA_193(.i_a(w_sum_128), .i_b(w_carry_165), .i_c(w_sum_166), .ow_sum(w_sum_193), .ow_carry(w_carry_193));
wire w_sum_194, w_carry_194;
math_adder_carry_save CSA_194(.i_a(w_sum_130), .i_b(w_carry_166), .i_c(w_sum_167), .ow_sum(w_sum_194), .ow_carry(w_carry_194));
wire w_sum_195, w_carry_195;
math_adder_carry_save CSA_195(.i_a(w_sum_132), .i_b(w_carry_167), .i_c(w_sum_168), .ow_sum(w_sum_195), .ow_carry(w_carry_195));
wire w_sum_196, w_carry_196;
math_adder_carry_save CSA_196(.i_a(w_sum_134), .i_b(w_carry_168), .i_c(w_sum_169), .ow_sum(w_sum_196), .ow_carry(w_carry_196));
wire w_sum_197, w_carry_197;
math_adder_carry_save CSA_197(.i_a(w_sum_136), .i_b(w_carry_169), .i_c(w_sum_170), .ow_sum(w_sum_197), .ow_carry(w_carry_197));
wire w_sum_198, w_carry_198;
math_adder_carry_save CSA_198(.i_a(w_sum_138), .i_b(w_carry_170), .i_c(w_sum_171), .ow_sum(w_sum_198), .ow_carry(w_carry_198));
wire w_sum_199, w_carry_199;
math_adder_carry_save CSA_199(.i_a(w_sum_140), .i_b(w_carry_171), .i_c(w_sum_172), .ow_sum(w_sum_199), .ow_carry(w_carry_199));
wire w_sum_200, w_carry_200;
math_adder_carry_save CSA_200(.i_a(w_sum_142), .i_b(w_carry_172), .i_c(w_sum_173), .ow_sum(w_sum_200), .ow_carry(w_carry_200));
wire w_sum_201, w_carry_201;
math_adder_carry_save CSA_201(.i_a(w_sum_144), .i_b(w_carry_173), .i_c(w_sum_174), .ow_sum(w_sum_201), .ow_carry(w_carry_201));
wire w_sum_202, w_carry_202;
math_adder_carry_save CSA_202(.i_a(w_sum_146), .i_b(w_carry_174), .i_c(w_sum_175), .ow_sum(w_sum_202), .ow_carry(w_carry_202));
wire w_sum_203, w_carry_203;
math_adder_carry_save CSA_203(.i_a(w_sum_148), .i_b(w_carry_175), .i_c(w_sum_176), .ow_sum(w_sum_203), .ow_carry(w_carry_203));
wire w_sum_204, w_carry_204;
math_adder_carry_save CSA_204(.i_a(w_sum_150), .i_b(w_carry_176), .i_c(w_sum_177), .ow_sum(w_sum_204), .ow_carry(w_carry_204));
wire w_sum_205, w_carry_205;
math_adder_carry_save CSA_205(.i_a(w_sum_152), .i_b(w_carry_177), .i_c(w_sum_178), .ow_sum(w_sum_205), .ow_carry(w_carry_205));
wire w_sum_206, w_carry_206;
math_adder_carry_save CSA_206(.i_a(w_sum_154), .i_b(w_carry_178), .i_c(w_sum_179), .ow_sum(w_sum_206), .ow_carry(w_carry_206));
wire w_sum_207, w_carry_207;
math_adder_carry_save CSA_207(.i_a(w_sum_155), .i_b(w_carry_179), .i_c(w_sum_180), .ow_sum(w_sum_207), .ow_carry(w_carry_207));
wire w_sum_208, w_carry_208;
math_adder_carry_save CSA_208(.i_a(w_carry_155), .i_b(w_carry_180), .i_c(w_sum_181), .ow_sum(w_sum_208), .ow_carry(w_carry_208));
wire w_sum_209, w_carry_209;
math_adder_carry_save CSA_209(.i_a(w_pp_14_15), .i_b(w_pp_15_14), .i_c(w_carry_181), .ow_sum(w_sum_209), .ow_carry(w_carry_209));

// Final addition stage
wire ow_sum_00, ow_carry_00;
assign ow_sum_00 = w_pp_00_00;
assign ow_carry_00 = 1'b0;
wire ow_sum_01, ow_carry_01;
math_adder_full FA_01(.i_a(w_pp_00_01), .i_b(w_pp_01_00), .i_c(ow_carry_00), .ow_sum(ow_sum_01), .ow_carry(ow_carry_01));
wire ow_sum_02, ow_carry_02;
math_adder_full FA_02(.i_a(w_pp_02_00), .i_b(w_sum_182), .i_c(ow_carry_01), .ow_sum(ow_sum_02), .ow_carry(ow_carry_02));
wire ow_sum_03, ow_carry_03;
math_adder_full FA_03(.i_a(w_carry_182), .i_b(w_sum_183), .i_c(ow_carry_02), .ow_sum(ow_sum_03), .ow_carry(ow_carry_03));
wire ow_sum_04, ow_carry_04;
math_adder_full FA_04(.i_a(w_carry_183), .i_b(w_sum_184), .i_c(ow_carry_03), .ow_sum(ow_sum_04), .ow_carry(ow_carry_04));
wire ow_sum_05, ow_carry_05;
math_adder_full FA_05(.i_a(w_carry_184), .i_b(w_sum_185), .i_c(ow_carry_04), .ow_sum(ow_sum_05), .ow_carry(ow_carry_05));
wire ow_sum_06, ow_carry_06;
math_adder_full FA_06(.i_a(w_carry_185), .i_b(w_sum_186), .i_c(ow_carry_05), .ow_sum(ow_sum_06), .ow_carry(ow_carry_06));
wire ow_sum_07, ow_carry_07;
math_adder_full FA_07(.i_a(w_carry_186), .i_b(w_sum_187), .i_c(ow_carry_06), .ow_sum(ow_sum_07), .ow_carry(ow_carry_07));
wire ow_sum_08, ow_carry_08;
math_adder_full FA_08(.i_a(w_carry_187), .i_b(w_sum_188), .i_c(ow_carry_07), .ow_sum(ow_sum_08), .ow_carry(ow_carry_08));
wire ow_sum_09, ow_carry_09;
math_adder_full FA_09(.i_a(w_carry_188), .i_b(w_sum_189), .i_c(ow_carry_08), .ow_sum(ow_sum_09), .ow_carry(ow_carry_09));
wire ow_sum_10, ow_carry_10;
math_adder_full FA_10(.i_a(w_carry_189), .i_b(w_sum_190), .i_c(ow_carry_09), .ow_sum(ow_sum_10), .ow_carry(ow_carry_10));
wire ow_sum_11, ow_carry_11;
math_adder_full FA_11(.i_a(w_carry_190), .i_b(w_sum_191), .i_c(ow_carry_10), .ow_sum(ow_sum_11), .ow_carry(ow_carry_11));
wire ow_sum_12, ow_carry_12;
math_adder_full FA_12(.i_a(w_carry_191), .i_b(w_sum_192), .i_c(ow_carry_11), .ow_sum(ow_sum_12), .ow_carry(ow_carry_12));
wire ow_sum_13, ow_carry_13;
math_adder_full FA_13(.i_a(w_carry_192), .i_b(w_sum_193), .i_c(ow_carry_12), .ow_sum(ow_sum_13), .ow_carry(ow_carry_13));
wire ow_sum_14, ow_carry_14;
math_adder_full FA_14(.i_a(w_carry_193), .i_b(w_sum_194), .i_c(ow_carry_13), .ow_sum(ow_sum_14), .ow_carry(ow_carry_14));
wire ow_sum_15, ow_carry_15;
math_adder_full FA_15(.i_a(w_carry_194), .i_b(w_sum_195), .i_c(ow_carry_14), .ow_sum(ow_sum_15), .ow_carry(ow_carry_15));
wire ow_sum_16, ow_carry_16;
math_adder_full FA_16(.i_a(w_carry_195), .i_b(w_sum_196), .i_c(ow_carry_15), .ow_sum(ow_sum_16), .ow_carry(ow_carry_16));
wire ow_sum_17, ow_carry_17;
math_adder_full FA_17(.i_a(w_carry_196), .i_b(w_sum_197), .i_c(ow_carry_16), .ow_sum(ow_sum_17), .ow_carry(ow_carry_17));
wire ow_sum_18, ow_carry_18;
math_adder_full FA_18(.i_a(w_carry_197), .i_b(w_sum_198), .i_c(ow_carry_17), .ow_sum(ow_sum_18), .ow_carry(ow_carry_18));
wire ow_sum_19, ow_carry_19;
math_adder_full FA_19(.i_a(w_carry_198), .i_b(w_sum_199), .i_c(ow_carry_18), .ow_sum(ow_sum_19), .ow_carry(ow_carry_19));
wire ow_sum_20, ow_carry_20;
math_adder_full FA_20(.i_a(w_carry_199), .i_b(w_sum_200), .i_c(ow_carry_19), .ow_sum(ow_sum_20), .ow_carry(ow_carry_20));
wire ow_sum_21, ow_carry_21;
math_adder_full FA_21(.i_a(w_carry_200), .i_b(w_sum_201), .i_c(ow_carry_20), .ow_sum(ow_sum_21), .ow_carry(ow_carry_21));
wire ow_sum_22, ow_carry_22;
math_adder_full FA_22(.i_a(w_carry_201), .i_b(w_sum_202), .i_c(ow_carry_21), .ow_sum(ow_sum_22), .ow_carry(ow_carry_22));
wire ow_sum_23, ow_carry_23;
math_adder_full FA_23(.i_a(w_carry_202), .i_b(w_sum_203), .i_c(ow_carry_22), .ow_sum(ow_sum_23), .ow_carry(ow_carry_23));
wire ow_sum_24, ow_carry_24;
math_adder_full FA_24(.i_a(w_carry_203), .i_b(w_sum_204), .i_c(ow_carry_23), .ow_sum(ow_sum_24), .ow_carry(ow_carry_24));
wire ow_sum_25, ow_carry_25;
math_adder_full FA_25(.i_a(w_carry_204), .i_b(w_sum_205), .i_c(ow_carry_24), .ow_sum(ow_sum_25), .ow_carry(ow_carry_25));
wire ow_sum_26, ow_carry_26;
math_adder_full FA_26(.i_a(w_carry_205), .i_b(w_sum_206), .i_c(ow_carry_25), .ow_sum(ow_sum_26), .ow_carry(ow_carry_26));
wire ow_sum_27, ow_carry_27;
math_adder_full FA_27(.i_a(w_carry_206), .i_b(w_sum_207), .i_c(ow_carry_26), .ow_sum(ow_sum_27), .ow_carry(ow_carry_27));
wire ow_sum_28, ow_carry_28;
math_adder_full FA_28(.i_a(w_carry_207), .i_b(w_sum_208), .i_c(ow_carry_27), .ow_sum(ow_sum_28), .ow_carry(ow_carry_28));
wire ow_sum_29, ow_carry_29;
math_adder_full FA_29(.i_a(w_carry_208), .i_b(w_sum_209), .i_c(ow_carry_28), .ow_sum(ow_sum_29), .ow_carry(ow_carry_29));
wire ow_sum_30, ow_carry_30;
math_adder_full FA_30(.i_a(w_pp_15_15), .i_b(w_carry_209), .i_c(ow_carry_29), .ow_sum(ow_sum_30), .ow_carry(ow_carry_30));
wire ow_sum_31, ow_carry_31;
assign ow_sum_31 = ow_carry_30;
assign ow_carry_31 = 1'b0;

// Final product assignment
assign ow_product[ 0] = ow_sum_00;
assign ow_product[ 1] = ow_sum_01;
assign ow_product[ 2] = ow_sum_02;
assign ow_product[ 3] = ow_sum_03;
assign ow_product[ 4] = ow_sum_04;
assign ow_product[ 5] = ow_sum_05;
assign ow_product[ 6] = ow_sum_06;
assign ow_product[ 7] = ow_sum_07;
assign ow_product[ 8] = ow_sum_08;
assign ow_product[ 9] = ow_sum_09;
assign ow_product[10] = ow_sum_10;
assign ow_product[11] = ow_sum_11;
assign ow_product[12] = ow_sum_12;
assign ow_product[13] = ow_sum_13;
assign ow_product[14] = ow_sum_14;
assign ow_product[15] = ow_sum_15;
assign ow_product[16] = ow_sum_16;
assign ow_product[17] = ow_sum_17;
assign ow_product[18] = ow_sum_18;
assign ow_product[19] = ow_sum_19;
assign ow_product[20] = ow_sum_20;
assign ow_product[21] = ow_sum_21;
assign ow_product[22] = ow_sum_22;
assign ow_product[23] = ow_sum_23;
assign ow_product[24] = ow_sum_24;
assign ow_product[25] = ow_sum_25;
assign ow_product[26] = ow_sum_26;
assign ow_product[27] = ow_sum_27;
assign ow_product[28] = ow_sum_28;
assign ow_product[29] = ow_sum_29;
assign ow_product[30] = ow_sum_30;
assign ow_product[31] = ow_sum_31;


    // Debug purposes
    // synopsys translate_off
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_dadda_tree_016);
    end
    // synopsys translate_on
        
endmodule : math_multiplier_dadda_tree_016
