`timescale 1ns / 1ps

module math_multiplier_dadda_tree_32 (
    input  [31:0] i_multiplier,
    input  [31:0] i_multiplicand,
    output [63:0] ow_product
);

// Partial products generation
wire w_pp_00_00 = i_multiplier[ 0] & i_multiplicand[ 0];
wire w_pp_00_01 = i_multiplier[ 0] & i_multiplicand[ 1];
wire w_pp_00_02 = i_multiplier[ 0] & i_multiplicand[ 2];
wire w_pp_00_03 = i_multiplier[ 0] & i_multiplicand[ 3];
wire w_pp_00_04 = i_multiplier[ 0] & i_multiplicand[ 4];
wire w_pp_00_05 = i_multiplier[ 0] & i_multiplicand[ 5];
wire w_pp_00_06 = i_multiplier[ 0] & i_multiplicand[ 6];
wire w_pp_00_07 = i_multiplier[ 0] & i_multiplicand[ 7];
wire w_pp_00_08 = i_multiplier[ 0] & i_multiplicand[ 8];
wire w_pp_00_09 = i_multiplier[ 0] & i_multiplicand[ 9];
wire w_pp_00_10 = i_multiplier[ 0] & i_multiplicand[10];
wire w_pp_00_11 = i_multiplier[ 0] & i_multiplicand[11];
wire w_pp_00_12 = i_multiplier[ 0] & i_multiplicand[12];
wire w_pp_00_13 = i_multiplier[ 0] & i_multiplicand[13];
wire w_pp_00_14 = i_multiplier[ 0] & i_multiplicand[14];
wire w_pp_00_15 = i_multiplier[ 0] & i_multiplicand[15];
wire w_pp_00_16 = i_multiplier[ 0] & i_multiplicand[16];
wire w_pp_00_17 = i_multiplier[ 0] & i_multiplicand[17];
wire w_pp_00_18 = i_multiplier[ 0] & i_multiplicand[18];
wire w_pp_00_19 = i_multiplier[ 0] & i_multiplicand[19];
wire w_pp_00_20 = i_multiplier[ 0] & i_multiplicand[20];
wire w_pp_00_21 = i_multiplier[ 0] & i_multiplicand[21];
wire w_pp_00_22 = i_multiplier[ 0] & i_multiplicand[22];
wire w_pp_00_23 = i_multiplier[ 0] & i_multiplicand[23];
wire w_pp_00_24 = i_multiplier[ 0] & i_multiplicand[24];
wire w_pp_00_25 = i_multiplier[ 0] & i_multiplicand[25];
wire w_pp_00_26 = i_multiplier[ 0] & i_multiplicand[26];
wire w_pp_00_27 = i_multiplier[ 0] & i_multiplicand[27];
wire w_pp_00_28 = i_multiplier[ 0] & i_multiplicand[28];
wire w_pp_00_29 = i_multiplier[ 0] & i_multiplicand[29];
wire w_pp_00_30 = i_multiplier[ 0] & i_multiplicand[30];
wire w_pp_00_31 = i_multiplier[ 0] & i_multiplicand[31];
wire w_pp_01_00 = i_multiplier[ 1] & i_multiplicand[ 0];
wire w_pp_01_01 = i_multiplier[ 1] & i_multiplicand[ 1];
wire w_pp_01_02 = i_multiplier[ 1] & i_multiplicand[ 2];
wire w_pp_01_03 = i_multiplier[ 1] & i_multiplicand[ 3];
wire w_pp_01_04 = i_multiplier[ 1] & i_multiplicand[ 4];
wire w_pp_01_05 = i_multiplier[ 1] & i_multiplicand[ 5];
wire w_pp_01_06 = i_multiplier[ 1] & i_multiplicand[ 6];
wire w_pp_01_07 = i_multiplier[ 1] & i_multiplicand[ 7];
wire w_pp_01_08 = i_multiplier[ 1] & i_multiplicand[ 8];
wire w_pp_01_09 = i_multiplier[ 1] & i_multiplicand[ 9];
wire w_pp_01_10 = i_multiplier[ 1] & i_multiplicand[10];
wire w_pp_01_11 = i_multiplier[ 1] & i_multiplicand[11];
wire w_pp_01_12 = i_multiplier[ 1] & i_multiplicand[12];
wire w_pp_01_13 = i_multiplier[ 1] & i_multiplicand[13];
wire w_pp_01_14 = i_multiplier[ 1] & i_multiplicand[14];
wire w_pp_01_15 = i_multiplier[ 1] & i_multiplicand[15];
wire w_pp_01_16 = i_multiplier[ 1] & i_multiplicand[16];
wire w_pp_01_17 = i_multiplier[ 1] & i_multiplicand[17];
wire w_pp_01_18 = i_multiplier[ 1] & i_multiplicand[18];
wire w_pp_01_19 = i_multiplier[ 1] & i_multiplicand[19];
wire w_pp_01_20 = i_multiplier[ 1] & i_multiplicand[20];
wire w_pp_01_21 = i_multiplier[ 1] & i_multiplicand[21];
wire w_pp_01_22 = i_multiplier[ 1] & i_multiplicand[22];
wire w_pp_01_23 = i_multiplier[ 1] & i_multiplicand[23];
wire w_pp_01_24 = i_multiplier[ 1] & i_multiplicand[24];
wire w_pp_01_25 = i_multiplier[ 1] & i_multiplicand[25];
wire w_pp_01_26 = i_multiplier[ 1] & i_multiplicand[26];
wire w_pp_01_27 = i_multiplier[ 1] & i_multiplicand[27];
wire w_pp_01_28 = i_multiplier[ 1] & i_multiplicand[28];
wire w_pp_01_29 = i_multiplier[ 1] & i_multiplicand[29];
wire w_pp_01_30 = i_multiplier[ 1] & i_multiplicand[30];
wire w_pp_01_31 = i_multiplier[ 1] & i_multiplicand[31];
wire w_pp_02_00 = i_multiplier[ 2] & i_multiplicand[ 0];
wire w_pp_02_01 = i_multiplier[ 2] & i_multiplicand[ 1];
wire w_pp_02_02 = i_multiplier[ 2] & i_multiplicand[ 2];
wire w_pp_02_03 = i_multiplier[ 2] & i_multiplicand[ 3];
wire w_pp_02_04 = i_multiplier[ 2] & i_multiplicand[ 4];
wire w_pp_02_05 = i_multiplier[ 2] & i_multiplicand[ 5];
wire w_pp_02_06 = i_multiplier[ 2] & i_multiplicand[ 6];
wire w_pp_02_07 = i_multiplier[ 2] & i_multiplicand[ 7];
wire w_pp_02_08 = i_multiplier[ 2] & i_multiplicand[ 8];
wire w_pp_02_09 = i_multiplier[ 2] & i_multiplicand[ 9];
wire w_pp_02_10 = i_multiplier[ 2] & i_multiplicand[10];
wire w_pp_02_11 = i_multiplier[ 2] & i_multiplicand[11];
wire w_pp_02_12 = i_multiplier[ 2] & i_multiplicand[12];
wire w_pp_02_13 = i_multiplier[ 2] & i_multiplicand[13];
wire w_pp_02_14 = i_multiplier[ 2] & i_multiplicand[14];
wire w_pp_02_15 = i_multiplier[ 2] & i_multiplicand[15];
wire w_pp_02_16 = i_multiplier[ 2] & i_multiplicand[16];
wire w_pp_02_17 = i_multiplier[ 2] & i_multiplicand[17];
wire w_pp_02_18 = i_multiplier[ 2] & i_multiplicand[18];
wire w_pp_02_19 = i_multiplier[ 2] & i_multiplicand[19];
wire w_pp_02_20 = i_multiplier[ 2] & i_multiplicand[20];
wire w_pp_02_21 = i_multiplier[ 2] & i_multiplicand[21];
wire w_pp_02_22 = i_multiplier[ 2] & i_multiplicand[22];
wire w_pp_02_23 = i_multiplier[ 2] & i_multiplicand[23];
wire w_pp_02_24 = i_multiplier[ 2] & i_multiplicand[24];
wire w_pp_02_25 = i_multiplier[ 2] & i_multiplicand[25];
wire w_pp_02_26 = i_multiplier[ 2] & i_multiplicand[26];
wire w_pp_02_27 = i_multiplier[ 2] & i_multiplicand[27];
wire w_pp_02_28 = i_multiplier[ 2] & i_multiplicand[28];
wire w_pp_02_29 = i_multiplier[ 2] & i_multiplicand[29];
wire w_pp_02_30 = i_multiplier[ 2] & i_multiplicand[30];
wire w_pp_02_31 = i_multiplier[ 2] & i_multiplicand[31];
wire w_pp_03_00 = i_multiplier[ 3] & i_multiplicand[ 0];
wire w_pp_03_01 = i_multiplier[ 3] & i_multiplicand[ 1];
wire w_pp_03_02 = i_multiplier[ 3] & i_multiplicand[ 2];
wire w_pp_03_03 = i_multiplier[ 3] & i_multiplicand[ 3];
wire w_pp_03_04 = i_multiplier[ 3] & i_multiplicand[ 4];
wire w_pp_03_05 = i_multiplier[ 3] & i_multiplicand[ 5];
wire w_pp_03_06 = i_multiplier[ 3] & i_multiplicand[ 6];
wire w_pp_03_07 = i_multiplier[ 3] & i_multiplicand[ 7];
wire w_pp_03_08 = i_multiplier[ 3] & i_multiplicand[ 8];
wire w_pp_03_09 = i_multiplier[ 3] & i_multiplicand[ 9];
wire w_pp_03_10 = i_multiplier[ 3] & i_multiplicand[10];
wire w_pp_03_11 = i_multiplier[ 3] & i_multiplicand[11];
wire w_pp_03_12 = i_multiplier[ 3] & i_multiplicand[12];
wire w_pp_03_13 = i_multiplier[ 3] & i_multiplicand[13];
wire w_pp_03_14 = i_multiplier[ 3] & i_multiplicand[14];
wire w_pp_03_15 = i_multiplier[ 3] & i_multiplicand[15];
wire w_pp_03_16 = i_multiplier[ 3] & i_multiplicand[16];
wire w_pp_03_17 = i_multiplier[ 3] & i_multiplicand[17];
wire w_pp_03_18 = i_multiplier[ 3] & i_multiplicand[18];
wire w_pp_03_19 = i_multiplier[ 3] & i_multiplicand[19];
wire w_pp_03_20 = i_multiplier[ 3] & i_multiplicand[20];
wire w_pp_03_21 = i_multiplier[ 3] & i_multiplicand[21];
wire w_pp_03_22 = i_multiplier[ 3] & i_multiplicand[22];
wire w_pp_03_23 = i_multiplier[ 3] & i_multiplicand[23];
wire w_pp_03_24 = i_multiplier[ 3] & i_multiplicand[24];
wire w_pp_03_25 = i_multiplier[ 3] & i_multiplicand[25];
wire w_pp_03_26 = i_multiplier[ 3] & i_multiplicand[26];
wire w_pp_03_27 = i_multiplier[ 3] & i_multiplicand[27];
wire w_pp_03_28 = i_multiplier[ 3] & i_multiplicand[28];
wire w_pp_03_29 = i_multiplier[ 3] & i_multiplicand[29];
wire w_pp_03_30 = i_multiplier[ 3] & i_multiplicand[30];
wire w_pp_03_31 = i_multiplier[ 3] & i_multiplicand[31];
wire w_pp_04_00 = i_multiplier[ 4] & i_multiplicand[ 0];
wire w_pp_04_01 = i_multiplier[ 4] & i_multiplicand[ 1];
wire w_pp_04_02 = i_multiplier[ 4] & i_multiplicand[ 2];
wire w_pp_04_03 = i_multiplier[ 4] & i_multiplicand[ 3];
wire w_pp_04_04 = i_multiplier[ 4] & i_multiplicand[ 4];
wire w_pp_04_05 = i_multiplier[ 4] & i_multiplicand[ 5];
wire w_pp_04_06 = i_multiplier[ 4] & i_multiplicand[ 6];
wire w_pp_04_07 = i_multiplier[ 4] & i_multiplicand[ 7];
wire w_pp_04_08 = i_multiplier[ 4] & i_multiplicand[ 8];
wire w_pp_04_09 = i_multiplier[ 4] & i_multiplicand[ 9];
wire w_pp_04_10 = i_multiplier[ 4] & i_multiplicand[10];
wire w_pp_04_11 = i_multiplier[ 4] & i_multiplicand[11];
wire w_pp_04_12 = i_multiplier[ 4] & i_multiplicand[12];
wire w_pp_04_13 = i_multiplier[ 4] & i_multiplicand[13];
wire w_pp_04_14 = i_multiplier[ 4] & i_multiplicand[14];
wire w_pp_04_15 = i_multiplier[ 4] & i_multiplicand[15];
wire w_pp_04_16 = i_multiplier[ 4] & i_multiplicand[16];
wire w_pp_04_17 = i_multiplier[ 4] & i_multiplicand[17];
wire w_pp_04_18 = i_multiplier[ 4] & i_multiplicand[18];
wire w_pp_04_19 = i_multiplier[ 4] & i_multiplicand[19];
wire w_pp_04_20 = i_multiplier[ 4] & i_multiplicand[20];
wire w_pp_04_21 = i_multiplier[ 4] & i_multiplicand[21];
wire w_pp_04_22 = i_multiplier[ 4] & i_multiplicand[22];
wire w_pp_04_23 = i_multiplier[ 4] & i_multiplicand[23];
wire w_pp_04_24 = i_multiplier[ 4] & i_multiplicand[24];
wire w_pp_04_25 = i_multiplier[ 4] & i_multiplicand[25];
wire w_pp_04_26 = i_multiplier[ 4] & i_multiplicand[26];
wire w_pp_04_27 = i_multiplier[ 4] & i_multiplicand[27];
wire w_pp_04_28 = i_multiplier[ 4] & i_multiplicand[28];
wire w_pp_04_29 = i_multiplier[ 4] & i_multiplicand[29];
wire w_pp_04_30 = i_multiplier[ 4] & i_multiplicand[30];
wire w_pp_04_31 = i_multiplier[ 4] & i_multiplicand[31];
wire w_pp_05_00 = i_multiplier[ 5] & i_multiplicand[ 0];
wire w_pp_05_01 = i_multiplier[ 5] & i_multiplicand[ 1];
wire w_pp_05_02 = i_multiplier[ 5] & i_multiplicand[ 2];
wire w_pp_05_03 = i_multiplier[ 5] & i_multiplicand[ 3];
wire w_pp_05_04 = i_multiplier[ 5] & i_multiplicand[ 4];
wire w_pp_05_05 = i_multiplier[ 5] & i_multiplicand[ 5];
wire w_pp_05_06 = i_multiplier[ 5] & i_multiplicand[ 6];
wire w_pp_05_07 = i_multiplier[ 5] & i_multiplicand[ 7];
wire w_pp_05_08 = i_multiplier[ 5] & i_multiplicand[ 8];
wire w_pp_05_09 = i_multiplier[ 5] & i_multiplicand[ 9];
wire w_pp_05_10 = i_multiplier[ 5] & i_multiplicand[10];
wire w_pp_05_11 = i_multiplier[ 5] & i_multiplicand[11];
wire w_pp_05_12 = i_multiplier[ 5] & i_multiplicand[12];
wire w_pp_05_13 = i_multiplier[ 5] & i_multiplicand[13];
wire w_pp_05_14 = i_multiplier[ 5] & i_multiplicand[14];
wire w_pp_05_15 = i_multiplier[ 5] & i_multiplicand[15];
wire w_pp_05_16 = i_multiplier[ 5] & i_multiplicand[16];
wire w_pp_05_17 = i_multiplier[ 5] & i_multiplicand[17];
wire w_pp_05_18 = i_multiplier[ 5] & i_multiplicand[18];
wire w_pp_05_19 = i_multiplier[ 5] & i_multiplicand[19];
wire w_pp_05_20 = i_multiplier[ 5] & i_multiplicand[20];
wire w_pp_05_21 = i_multiplier[ 5] & i_multiplicand[21];
wire w_pp_05_22 = i_multiplier[ 5] & i_multiplicand[22];
wire w_pp_05_23 = i_multiplier[ 5] & i_multiplicand[23];
wire w_pp_05_24 = i_multiplier[ 5] & i_multiplicand[24];
wire w_pp_05_25 = i_multiplier[ 5] & i_multiplicand[25];
wire w_pp_05_26 = i_multiplier[ 5] & i_multiplicand[26];
wire w_pp_05_27 = i_multiplier[ 5] & i_multiplicand[27];
wire w_pp_05_28 = i_multiplier[ 5] & i_multiplicand[28];
wire w_pp_05_29 = i_multiplier[ 5] & i_multiplicand[29];
wire w_pp_05_30 = i_multiplier[ 5] & i_multiplicand[30];
wire w_pp_05_31 = i_multiplier[ 5] & i_multiplicand[31];
wire w_pp_06_00 = i_multiplier[ 6] & i_multiplicand[ 0];
wire w_pp_06_01 = i_multiplier[ 6] & i_multiplicand[ 1];
wire w_pp_06_02 = i_multiplier[ 6] & i_multiplicand[ 2];
wire w_pp_06_03 = i_multiplier[ 6] & i_multiplicand[ 3];
wire w_pp_06_04 = i_multiplier[ 6] & i_multiplicand[ 4];
wire w_pp_06_05 = i_multiplier[ 6] & i_multiplicand[ 5];
wire w_pp_06_06 = i_multiplier[ 6] & i_multiplicand[ 6];
wire w_pp_06_07 = i_multiplier[ 6] & i_multiplicand[ 7];
wire w_pp_06_08 = i_multiplier[ 6] & i_multiplicand[ 8];
wire w_pp_06_09 = i_multiplier[ 6] & i_multiplicand[ 9];
wire w_pp_06_10 = i_multiplier[ 6] & i_multiplicand[10];
wire w_pp_06_11 = i_multiplier[ 6] & i_multiplicand[11];
wire w_pp_06_12 = i_multiplier[ 6] & i_multiplicand[12];
wire w_pp_06_13 = i_multiplier[ 6] & i_multiplicand[13];
wire w_pp_06_14 = i_multiplier[ 6] & i_multiplicand[14];
wire w_pp_06_15 = i_multiplier[ 6] & i_multiplicand[15];
wire w_pp_06_16 = i_multiplier[ 6] & i_multiplicand[16];
wire w_pp_06_17 = i_multiplier[ 6] & i_multiplicand[17];
wire w_pp_06_18 = i_multiplier[ 6] & i_multiplicand[18];
wire w_pp_06_19 = i_multiplier[ 6] & i_multiplicand[19];
wire w_pp_06_20 = i_multiplier[ 6] & i_multiplicand[20];
wire w_pp_06_21 = i_multiplier[ 6] & i_multiplicand[21];
wire w_pp_06_22 = i_multiplier[ 6] & i_multiplicand[22];
wire w_pp_06_23 = i_multiplier[ 6] & i_multiplicand[23];
wire w_pp_06_24 = i_multiplier[ 6] & i_multiplicand[24];
wire w_pp_06_25 = i_multiplier[ 6] & i_multiplicand[25];
wire w_pp_06_26 = i_multiplier[ 6] & i_multiplicand[26];
wire w_pp_06_27 = i_multiplier[ 6] & i_multiplicand[27];
wire w_pp_06_28 = i_multiplier[ 6] & i_multiplicand[28];
wire w_pp_06_29 = i_multiplier[ 6] & i_multiplicand[29];
wire w_pp_06_30 = i_multiplier[ 6] & i_multiplicand[30];
wire w_pp_06_31 = i_multiplier[ 6] & i_multiplicand[31];
wire w_pp_07_00 = i_multiplier[ 7] & i_multiplicand[ 0];
wire w_pp_07_01 = i_multiplier[ 7] & i_multiplicand[ 1];
wire w_pp_07_02 = i_multiplier[ 7] & i_multiplicand[ 2];
wire w_pp_07_03 = i_multiplier[ 7] & i_multiplicand[ 3];
wire w_pp_07_04 = i_multiplier[ 7] & i_multiplicand[ 4];
wire w_pp_07_05 = i_multiplier[ 7] & i_multiplicand[ 5];
wire w_pp_07_06 = i_multiplier[ 7] & i_multiplicand[ 6];
wire w_pp_07_07 = i_multiplier[ 7] & i_multiplicand[ 7];
wire w_pp_07_08 = i_multiplier[ 7] & i_multiplicand[ 8];
wire w_pp_07_09 = i_multiplier[ 7] & i_multiplicand[ 9];
wire w_pp_07_10 = i_multiplier[ 7] & i_multiplicand[10];
wire w_pp_07_11 = i_multiplier[ 7] & i_multiplicand[11];
wire w_pp_07_12 = i_multiplier[ 7] & i_multiplicand[12];
wire w_pp_07_13 = i_multiplier[ 7] & i_multiplicand[13];
wire w_pp_07_14 = i_multiplier[ 7] & i_multiplicand[14];
wire w_pp_07_15 = i_multiplier[ 7] & i_multiplicand[15];
wire w_pp_07_16 = i_multiplier[ 7] & i_multiplicand[16];
wire w_pp_07_17 = i_multiplier[ 7] & i_multiplicand[17];
wire w_pp_07_18 = i_multiplier[ 7] & i_multiplicand[18];
wire w_pp_07_19 = i_multiplier[ 7] & i_multiplicand[19];
wire w_pp_07_20 = i_multiplier[ 7] & i_multiplicand[20];
wire w_pp_07_21 = i_multiplier[ 7] & i_multiplicand[21];
wire w_pp_07_22 = i_multiplier[ 7] & i_multiplicand[22];
wire w_pp_07_23 = i_multiplier[ 7] & i_multiplicand[23];
wire w_pp_07_24 = i_multiplier[ 7] & i_multiplicand[24];
wire w_pp_07_25 = i_multiplier[ 7] & i_multiplicand[25];
wire w_pp_07_26 = i_multiplier[ 7] & i_multiplicand[26];
wire w_pp_07_27 = i_multiplier[ 7] & i_multiplicand[27];
wire w_pp_07_28 = i_multiplier[ 7] & i_multiplicand[28];
wire w_pp_07_29 = i_multiplier[ 7] & i_multiplicand[29];
wire w_pp_07_30 = i_multiplier[ 7] & i_multiplicand[30];
wire w_pp_07_31 = i_multiplier[ 7] & i_multiplicand[31];
wire w_pp_08_00 = i_multiplier[ 8] & i_multiplicand[ 0];
wire w_pp_08_01 = i_multiplier[ 8] & i_multiplicand[ 1];
wire w_pp_08_02 = i_multiplier[ 8] & i_multiplicand[ 2];
wire w_pp_08_03 = i_multiplier[ 8] & i_multiplicand[ 3];
wire w_pp_08_04 = i_multiplier[ 8] & i_multiplicand[ 4];
wire w_pp_08_05 = i_multiplier[ 8] & i_multiplicand[ 5];
wire w_pp_08_06 = i_multiplier[ 8] & i_multiplicand[ 6];
wire w_pp_08_07 = i_multiplier[ 8] & i_multiplicand[ 7];
wire w_pp_08_08 = i_multiplier[ 8] & i_multiplicand[ 8];
wire w_pp_08_09 = i_multiplier[ 8] & i_multiplicand[ 9];
wire w_pp_08_10 = i_multiplier[ 8] & i_multiplicand[10];
wire w_pp_08_11 = i_multiplier[ 8] & i_multiplicand[11];
wire w_pp_08_12 = i_multiplier[ 8] & i_multiplicand[12];
wire w_pp_08_13 = i_multiplier[ 8] & i_multiplicand[13];
wire w_pp_08_14 = i_multiplier[ 8] & i_multiplicand[14];
wire w_pp_08_15 = i_multiplier[ 8] & i_multiplicand[15];
wire w_pp_08_16 = i_multiplier[ 8] & i_multiplicand[16];
wire w_pp_08_17 = i_multiplier[ 8] & i_multiplicand[17];
wire w_pp_08_18 = i_multiplier[ 8] & i_multiplicand[18];
wire w_pp_08_19 = i_multiplier[ 8] & i_multiplicand[19];
wire w_pp_08_20 = i_multiplier[ 8] & i_multiplicand[20];
wire w_pp_08_21 = i_multiplier[ 8] & i_multiplicand[21];
wire w_pp_08_22 = i_multiplier[ 8] & i_multiplicand[22];
wire w_pp_08_23 = i_multiplier[ 8] & i_multiplicand[23];
wire w_pp_08_24 = i_multiplier[ 8] & i_multiplicand[24];
wire w_pp_08_25 = i_multiplier[ 8] & i_multiplicand[25];
wire w_pp_08_26 = i_multiplier[ 8] & i_multiplicand[26];
wire w_pp_08_27 = i_multiplier[ 8] & i_multiplicand[27];
wire w_pp_08_28 = i_multiplier[ 8] & i_multiplicand[28];
wire w_pp_08_29 = i_multiplier[ 8] & i_multiplicand[29];
wire w_pp_08_30 = i_multiplier[ 8] & i_multiplicand[30];
wire w_pp_08_31 = i_multiplier[ 8] & i_multiplicand[31];
wire w_pp_09_00 = i_multiplier[ 9] & i_multiplicand[ 0];
wire w_pp_09_01 = i_multiplier[ 9] & i_multiplicand[ 1];
wire w_pp_09_02 = i_multiplier[ 9] & i_multiplicand[ 2];
wire w_pp_09_03 = i_multiplier[ 9] & i_multiplicand[ 3];
wire w_pp_09_04 = i_multiplier[ 9] & i_multiplicand[ 4];
wire w_pp_09_05 = i_multiplier[ 9] & i_multiplicand[ 5];
wire w_pp_09_06 = i_multiplier[ 9] & i_multiplicand[ 6];
wire w_pp_09_07 = i_multiplier[ 9] & i_multiplicand[ 7];
wire w_pp_09_08 = i_multiplier[ 9] & i_multiplicand[ 8];
wire w_pp_09_09 = i_multiplier[ 9] & i_multiplicand[ 9];
wire w_pp_09_10 = i_multiplier[ 9] & i_multiplicand[10];
wire w_pp_09_11 = i_multiplier[ 9] & i_multiplicand[11];
wire w_pp_09_12 = i_multiplier[ 9] & i_multiplicand[12];
wire w_pp_09_13 = i_multiplier[ 9] & i_multiplicand[13];
wire w_pp_09_14 = i_multiplier[ 9] & i_multiplicand[14];
wire w_pp_09_15 = i_multiplier[ 9] & i_multiplicand[15];
wire w_pp_09_16 = i_multiplier[ 9] & i_multiplicand[16];
wire w_pp_09_17 = i_multiplier[ 9] & i_multiplicand[17];
wire w_pp_09_18 = i_multiplier[ 9] & i_multiplicand[18];
wire w_pp_09_19 = i_multiplier[ 9] & i_multiplicand[19];
wire w_pp_09_20 = i_multiplier[ 9] & i_multiplicand[20];
wire w_pp_09_21 = i_multiplier[ 9] & i_multiplicand[21];
wire w_pp_09_22 = i_multiplier[ 9] & i_multiplicand[22];
wire w_pp_09_23 = i_multiplier[ 9] & i_multiplicand[23];
wire w_pp_09_24 = i_multiplier[ 9] & i_multiplicand[24];
wire w_pp_09_25 = i_multiplier[ 9] & i_multiplicand[25];
wire w_pp_09_26 = i_multiplier[ 9] & i_multiplicand[26];
wire w_pp_09_27 = i_multiplier[ 9] & i_multiplicand[27];
wire w_pp_09_28 = i_multiplier[ 9] & i_multiplicand[28];
wire w_pp_09_29 = i_multiplier[ 9] & i_multiplicand[29];
wire w_pp_09_30 = i_multiplier[ 9] & i_multiplicand[30];
wire w_pp_09_31 = i_multiplier[ 9] & i_multiplicand[31];
wire w_pp_10_00 = i_multiplier[10] & i_multiplicand[ 0];
wire w_pp_10_01 = i_multiplier[10] & i_multiplicand[ 1];
wire w_pp_10_02 = i_multiplier[10] & i_multiplicand[ 2];
wire w_pp_10_03 = i_multiplier[10] & i_multiplicand[ 3];
wire w_pp_10_04 = i_multiplier[10] & i_multiplicand[ 4];
wire w_pp_10_05 = i_multiplier[10] & i_multiplicand[ 5];
wire w_pp_10_06 = i_multiplier[10] & i_multiplicand[ 6];
wire w_pp_10_07 = i_multiplier[10] & i_multiplicand[ 7];
wire w_pp_10_08 = i_multiplier[10] & i_multiplicand[ 8];
wire w_pp_10_09 = i_multiplier[10] & i_multiplicand[ 9];
wire w_pp_10_10 = i_multiplier[10] & i_multiplicand[10];
wire w_pp_10_11 = i_multiplier[10] & i_multiplicand[11];
wire w_pp_10_12 = i_multiplier[10] & i_multiplicand[12];
wire w_pp_10_13 = i_multiplier[10] & i_multiplicand[13];
wire w_pp_10_14 = i_multiplier[10] & i_multiplicand[14];
wire w_pp_10_15 = i_multiplier[10] & i_multiplicand[15];
wire w_pp_10_16 = i_multiplier[10] & i_multiplicand[16];
wire w_pp_10_17 = i_multiplier[10] & i_multiplicand[17];
wire w_pp_10_18 = i_multiplier[10] & i_multiplicand[18];
wire w_pp_10_19 = i_multiplier[10] & i_multiplicand[19];
wire w_pp_10_20 = i_multiplier[10] & i_multiplicand[20];
wire w_pp_10_21 = i_multiplier[10] & i_multiplicand[21];
wire w_pp_10_22 = i_multiplier[10] & i_multiplicand[22];
wire w_pp_10_23 = i_multiplier[10] & i_multiplicand[23];
wire w_pp_10_24 = i_multiplier[10] & i_multiplicand[24];
wire w_pp_10_25 = i_multiplier[10] & i_multiplicand[25];
wire w_pp_10_26 = i_multiplier[10] & i_multiplicand[26];
wire w_pp_10_27 = i_multiplier[10] & i_multiplicand[27];
wire w_pp_10_28 = i_multiplier[10] & i_multiplicand[28];
wire w_pp_10_29 = i_multiplier[10] & i_multiplicand[29];
wire w_pp_10_30 = i_multiplier[10] & i_multiplicand[30];
wire w_pp_10_31 = i_multiplier[10] & i_multiplicand[31];
wire w_pp_11_00 = i_multiplier[11] & i_multiplicand[ 0];
wire w_pp_11_01 = i_multiplier[11] & i_multiplicand[ 1];
wire w_pp_11_02 = i_multiplier[11] & i_multiplicand[ 2];
wire w_pp_11_03 = i_multiplier[11] & i_multiplicand[ 3];
wire w_pp_11_04 = i_multiplier[11] & i_multiplicand[ 4];
wire w_pp_11_05 = i_multiplier[11] & i_multiplicand[ 5];
wire w_pp_11_06 = i_multiplier[11] & i_multiplicand[ 6];
wire w_pp_11_07 = i_multiplier[11] & i_multiplicand[ 7];
wire w_pp_11_08 = i_multiplier[11] & i_multiplicand[ 8];
wire w_pp_11_09 = i_multiplier[11] & i_multiplicand[ 9];
wire w_pp_11_10 = i_multiplier[11] & i_multiplicand[10];
wire w_pp_11_11 = i_multiplier[11] & i_multiplicand[11];
wire w_pp_11_12 = i_multiplier[11] & i_multiplicand[12];
wire w_pp_11_13 = i_multiplier[11] & i_multiplicand[13];
wire w_pp_11_14 = i_multiplier[11] & i_multiplicand[14];
wire w_pp_11_15 = i_multiplier[11] & i_multiplicand[15];
wire w_pp_11_16 = i_multiplier[11] & i_multiplicand[16];
wire w_pp_11_17 = i_multiplier[11] & i_multiplicand[17];
wire w_pp_11_18 = i_multiplier[11] & i_multiplicand[18];
wire w_pp_11_19 = i_multiplier[11] & i_multiplicand[19];
wire w_pp_11_20 = i_multiplier[11] & i_multiplicand[20];
wire w_pp_11_21 = i_multiplier[11] & i_multiplicand[21];
wire w_pp_11_22 = i_multiplier[11] & i_multiplicand[22];
wire w_pp_11_23 = i_multiplier[11] & i_multiplicand[23];
wire w_pp_11_24 = i_multiplier[11] & i_multiplicand[24];
wire w_pp_11_25 = i_multiplier[11] & i_multiplicand[25];
wire w_pp_11_26 = i_multiplier[11] & i_multiplicand[26];
wire w_pp_11_27 = i_multiplier[11] & i_multiplicand[27];
wire w_pp_11_28 = i_multiplier[11] & i_multiplicand[28];
wire w_pp_11_29 = i_multiplier[11] & i_multiplicand[29];
wire w_pp_11_30 = i_multiplier[11] & i_multiplicand[30];
wire w_pp_11_31 = i_multiplier[11] & i_multiplicand[31];
wire w_pp_12_00 = i_multiplier[12] & i_multiplicand[ 0];
wire w_pp_12_01 = i_multiplier[12] & i_multiplicand[ 1];
wire w_pp_12_02 = i_multiplier[12] & i_multiplicand[ 2];
wire w_pp_12_03 = i_multiplier[12] & i_multiplicand[ 3];
wire w_pp_12_04 = i_multiplier[12] & i_multiplicand[ 4];
wire w_pp_12_05 = i_multiplier[12] & i_multiplicand[ 5];
wire w_pp_12_06 = i_multiplier[12] & i_multiplicand[ 6];
wire w_pp_12_07 = i_multiplier[12] & i_multiplicand[ 7];
wire w_pp_12_08 = i_multiplier[12] & i_multiplicand[ 8];
wire w_pp_12_09 = i_multiplier[12] & i_multiplicand[ 9];
wire w_pp_12_10 = i_multiplier[12] & i_multiplicand[10];
wire w_pp_12_11 = i_multiplier[12] & i_multiplicand[11];
wire w_pp_12_12 = i_multiplier[12] & i_multiplicand[12];
wire w_pp_12_13 = i_multiplier[12] & i_multiplicand[13];
wire w_pp_12_14 = i_multiplier[12] & i_multiplicand[14];
wire w_pp_12_15 = i_multiplier[12] & i_multiplicand[15];
wire w_pp_12_16 = i_multiplier[12] & i_multiplicand[16];
wire w_pp_12_17 = i_multiplier[12] & i_multiplicand[17];
wire w_pp_12_18 = i_multiplier[12] & i_multiplicand[18];
wire w_pp_12_19 = i_multiplier[12] & i_multiplicand[19];
wire w_pp_12_20 = i_multiplier[12] & i_multiplicand[20];
wire w_pp_12_21 = i_multiplier[12] & i_multiplicand[21];
wire w_pp_12_22 = i_multiplier[12] & i_multiplicand[22];
wire w_pp_12_23 = i_multiplier[12] & i_multiplicand[23];
wire w_pp_12_24 = i_multiplier[12] & i_multiplicand[24];
wire w_pp_12_25 = i_multiplier[12] & i_multiplicand[25];
wire w_pp_12_26 = i_multiplier[12] & i_multiplicand[26];
wire w_pp_12_27 = i_multiplier[12] & i_multiplicand[27];
wire w_pp_12_28 = i_multiplier[12] & i_multiplicand[28];
wire w_pp_12_29 = i_multiplier[12] & i_multiplicand[29];
wire w_pp_12_30 = i_multiplier[12] & i_multiplicand[30];
wire w_pp_12_31 = i_multiplier[12] & i_multiplicand[31];
wire w_pp_13_00 = i_multiplier[13] & i_multiplicand[ 0];
wire w_pp_13_01 = i_multiplier[13] & i_multiplicand[ 1];
wire w_pp_13_02 = i_multiplier[13] & i_multiplicand[ 2];
wire w_pp_13_03 = i_multiplier[13] & i_multiplicand[ 3];
wire w_pp_13_04 = i_multiplier[13] & i_multiplicand[ 4];
wire w_pp_13_05 = i_multiplier[13] & i_multiplicand[ 5];
wire w_pp_13_06 = i_multiplier[13] & i_multiplicand[ 6];
wire w_pp_13_07 = i_multiplier[13] & i_multiplicand[ 7];
wire w_pp_13_08 = i_multiplier[13] & i_multiplicand[ 8];
wire w_pp_13_09 = i_multiplier[13] & i_multiplicand[ 9];
wire w_pp_13_10 = i_multiplier[13] & i_multiplicand[10];
wire w_pp_13_11 = i_multiplier[13] & i_multiplicand[11];
wire w_pp_13_12 = i_multiplier[13] & i_multiplicand[12];
wire w_pp_13_13 = i_multiplier[13] & i_multiplicand[13];
wire w_pp_13_14 = i_multiplier[13] & i_multiplicand[14];
wire w_pp_13_15 = i_multiplier[13] & i_multiplicand[15];
wire w_pp_13_16 = i_multiplier[13] & i_multiplicand[16];
wire w_pp_13_17 = i_multiplier[13] & i_multiplicand[17];
wire w_pp_13_18 = i_multiplier[13] & i_multiplicand[18];
wire w_pp_13_19 = i_multiplier[13] & i_multiplicand[19];
wire w_pp_13_20 = i_multiplier[13] & i_multiplicand[20];
wire w_pp_13_21 = i_multiplier[13] & i_multiplicand[21];
wire w_pp_13_22 = i_multiplier[13] & i_multiplicand[22];
wire w_pp_13_23 = i_multiplier[13] & i_multiplicand[23];
wire w_pp_13_24 = i_multiplier[13] & i_multiplicand[24];
wire w_pp_13_25 = i_multiplier[13] & i_multiplicand[25];
wire w_pp_13_26 = i_multiplier[13] & i_multiplicand[26];
wire w_pp_13_27 = i_multiplier[13] & i_multiplicand[27];
wire w_pp_13_28 = i_multiplier[13] & i_multiplicand[28];
wire w_pp_13_29 = i_multiplier[13] & i_multiplicand[29];
wire w_pp_13_30 = i_multiplier[13] & i_multiplicand[30];
wire w_pp_13_31 = i_multiplier[13] & i_multiplicand[31];
wire w_pp_14_00 = i_multiplier[14] & i_multiplicand[ 0];
wire w_pp_14_01 = i_multiplier[14] & i_multiplicand[ 1];
wire w_pp_14_02 = i_multiplier[14] & i_multiplicand[ 2];
wire w_pp_14_03 = i_multiplier[14] & i_multiplicand[ 3];
wire w_pp_14_04 = i_multiplier[14] & i_multiplicand[ 4];
wire w_pp_14_05 = i_multiplier[14] & i_multiplicand[ 5];
wire w_pp_14_06 = i_multiplier[14] & i_multiplicand[ 6];
wire w_pp_14_07 = i_multiplier[14] & i_multiplicand[ 7];
wire w_pp_14_08 = i_multiplier[14] & i_multiplicand[ 8];
wire w_pp_14_09 = i_multiplier[14] & i_multiplicand[ 9];
wire w_pp_14_10 = i_multiplier[14] & i_multiplicand[10];
wire w_pp_14_11 = i_multiplier[14] & i_multiplicand[11];
wire w_pp_14_12 = i_multiplier[14] & i_multiplicand[12];
wire w_pp_14_13 = i_multiplier[14] & i_multiplicand[13];
wire w_pp_14_14 = i_multiplier[14] & i_multiplicand[14];
wire w_pp_14_15 = i_multiplier[14] & i_multiplicand[15];
wire w_pp_14_16 = i_multiplier[14] & i_multiplicand[16];
wire w_pp_14_17 = i_multiplier[14] & i_multiplicand[17];
wire w_pp_14_18 = i_multiplier[14] & i_multiplicand[18];
wire w_pp_14_19 = i_multiplier[14] & i_multiplicand[19];
wire w_pp_14_20 = i_multiplier[14] & i_multiplicand[20];
wire w_pp_14_21 = i_multiplier[14] & i_multiplicand[21];
wire w_pp_14_22 = i_multiplier[14] & i_multiplicand[22];
wire w_pp_14_23 = i_multiplier[14] & i_multiplicand[23];
wire w_pp_14_24 = i_multiplier[14] & i_multiplicand[24];
wire w_pp_14_25 = i_multiplier[14] & i_multiplicand[25];
wire w_pp_14_26 = i_multiplier[14] & i_multiplicand[26];
wire w_pp_14_27 = i_multiplier[14] & i_multiplicand[27];
wire w_pp_14_28 = i_multiplier[14] & i_multiplicand[28];
wire w_pp_14_29 = i_multiplier[14] & i_multiplicand[29];
wire w_pp_14_30 = i_multiplier[14] & i_multiplicand[30];
wire w_pp_14_31 = i_multiplier[14] & i_multiplicand[31];
wire w_pp_15_00 = i_multiplier[15] & i_multiplicand[ 0];
wire w_pp_15_01 = i_multiplier[15] & i_multiplicand[ 1];
wire w_pp_15_02 = i_multiplier[15] & i_multiplicand[ 2];
wire w_pp_15_03 = i_multiplier[15] & i_multiplicand[ 3];
wire w_pp_15_04 = i_multiplier[15] & i_multiplicand[ 4];
wire w_pp_15_05 = i_multiplier[15] & i_multiplicand[ 5];
wire w_pp_15_06 = i_multiplier[15] & i_multiplicand[ 6];
wire w_pp_15_07 = i_multiplier[15] & i_multiplicand[ 7];
wire w_pp_15_08 = i_multiplier[15] & i_multiplicand[ 8];
wire w_pp_15_09 = i_multiplier[15] & i_multiplicand[ 9];
wire w_pp_15_10 = i_multiplier[15] & i_multiplicand[10];
wire w_pp_15_11 = i_multiplier[15] & i_multiplicand[11];
wire w_pp_15_12 = i_multiplier[15] & i_multiplicand[12];
wire w_pp_15_13 = i_multiplier[15] & i_multiplicand[13];
wire w_pp_15_14 = i_multiplier[15] & i_multiplicand[14];
wire w_pp_15_15 = i_multiplier[15] & i_multiplicand[15];
wire w_pp_15_16 = i_multiplier[15] & i_multiplicand[16];
wire w_pp_15_17 = i_multiplier[15] & i_multiplicand[17];
wire w_pp_15_18 = i_multiplier[15] & i_multiplicand[18];
wire w_pp_15_19 = i_multiplier[15] & i_multiplicand[19];
wire w_pp_15_20 = i_multiplier[15] & i_multiplicand[20];
wire w_pp_15_21 = i_multiplier[15] & i_multiplicand[21];
wire w_pp_15_22 = i_multiplier[15] & i_multiplicand[22];
wire w_pp_15_23 = i_multiplier[15] & i_multiplicand[23];
wire w_pp_15_24 = i_multiplier[15] & i_multiplicand[24];
wire w_pp_15_25 = i_multiplier[15] & i_multiplicand[25];
wire w_pp_15_26 = i_multiplier[15] & i_multiplicand[26];
wire w_pp_15_27 = i_multiplier[15] & i_multiplicand[27];
wire w_pp_15_28 = i_multiplier[15] & i_multiplicand[28];
wire w_pp_15_29 = i_multiplier[15] & i_multiplicand[29];
wire w_pp_15_30 = i_multiplier[15] & i_multiplicand[30];
wire w_pp_15_31 = i_multiplier[15] & i_multiplicand[31];
wire w_pp_16_00 = i_multiplier[16] & i_multiplicand[ 0];
wire w_pp_16_01 = i_multiplier[16] & i_multiplicand[ 1];
wire w_pp_16_02 = i_multiplier[16] & i_multiplicand[ 2];
wire w_pp_16_03 = i_multiplier[16] & i_multiplicand[ 3];
wire w_pp_16_04 = i_multiplier[16] & i_multiplicand[ 4];
wire w_pp_16_05 = i_multiplier[16] & i_multiplicand[ 5];
wire w_pp_16_06 = i_multiplier[16] & i_multiplicand[ 6];
wire w_pp_16_07 = i_multiplier[16] & i_multiplicand[ 7];
wire w_pp_16_08 = i_multiplier[16] & i_multiplicand[ 8];
wire w_pp_16_09 = i_multiplier[16] & i_multiplicand[ 9];
wire w_pp_16_10 = i_multiplier[16] & i_multiplicand[10];
wire w_pp_16_11 = i_multiplier[16] & i_multiplicand[11];
wire w_pp_16_12 = i_multiplier[16] & i_multiplicand[12];
wire w_pp_16_13 = i_multiplier[16] & i_multiplicand[13];
wire w_pp_16_14 = i_multiplier[16] & i_multiplicand[14];
wire w_pp_16_15 = i_multiplier[16] & i_multiplicand[15];
wire w_pp_16_16 = i_multiplier[16] & i_multiplicand[16];
wire w_pp_16_17 = i_multiplier[16] & i_multiplicand[17];
wire w_pp_16_18 = i_multiplier[16] & i_multiplicand[18];
wire w_pp_16_19 = i_multiplier[16] & i_multiplicand[19];
wire w_pp_16_20 = i_multiplier[16] & i_multiplicand[20];
wire w_pp_16_21 = i_multiplier[16] & i_multiplicand[21];
wire w_pp_16_22 = i_multiplier[16] & i_multiplicand[22];
wire w_pp_16_23 = i_multiplier[16] & i_multiplicand[23];
wire w_pp_16_24 = i_multiplier[16] & i_multiplicand[24];
wire w_pp_16_25 = i_multiplier[16] & i_multiplicand[25];
wire w_pp_16_26 = i_multiplier[16] & i_multiplicand[26];
wire w_pp_16_27 = i_multiplier[16] & i_multiplicand[27];
wire w_pp_16_28 = i_multiplier[16] & i_multiplicand[28];
wire w_pp_16_29 = i_multiplier[16] & i_multiplicand[29];
wire w_pp_16_30 = i_multiplier[16] & i_multiplicand[30];
wire w_pp_16_31 = i_multiplier[16] & i_multiplicand[31];
wire w_pp_17_00 = i_multiplier[17] & i_multiplicand[ 0];
wire w_pp_17_01 = i_multiplier[17] & i_multiplicand[ 1];
wire w_pp_17_02 = i_multiplier[17] & i_multiplicand[ 2];
wire w_pp_17_03 = i_multiplier[17] & i_multiplicand[ 3];
wire w_pp_17_04 = i_multiplier[17] & i_multiplicand[ 4];
wire w_pp_17_05 = i_multiplier[17] & i_multiplicand[ 5];
wire w_pp_17_06 = i_multiplier[17] & i_multiplicand[ 6];
wire w_pp_17_07 = i_multiplier[17] & i_multiplicand[ 7];
wire w_pp_17_08 = i_multiplier[17] & i_multiplicand[ 8];
wire w_pp_17_09 = i_multiplier[17] & i_multiplicand[ 9];
wire w_pp_17_10 = i_multiplier[17] & i_multiplicand[10];
wire w_pp_17_11 = i_multiplier[17] & i_multiplicand[11];
wire w_pp_17_12 = i_multiplier[17] & i_multiplicand[12];
wire w_pp_17_13 = i_multiplier[17] & i_multiplicand[13];
wire w_pp_17_14 = i_multiplier[17] & i_multiplicand[14];
wire w_pp_17_15 = i_multiplier[17] & i_multiplicand[15];
wire w_pp_17_16 = i_multiplier[17] & i_multiplicand[16];
wire w_pp_17_17 = i_multiplier[17] & i_multiplicand[17];
wire w_pp_17_18 = i_multiplier[17] & i_multiplicand[18];
wire w_pp_17_19 = i_multiplier[17] & i_multiplicand[19];
wire w_pp_17_20 = i_multiplier[17] & i_multiplicand[20];
wire w_pp_17_21 = i_multiplier[17] & i_multiplicand[21];
wire w_pp_17_22 = i_multiplier[17] & i_multiplicand[22];
wire w_pp_17_23 = i_multiplier[17] & i_multiplicand[23];
wire w_pp_17_24 = i_multiplier[17] & i_multiplicand[24];
wire w_pp_17_25 = i_multiplier[17] & i_multiplicand[25];
wire w_pp_17_26 = i_multiplier[17] & i_multiplicand[26];
wire w_pp_17_27 = i_multiplier[17] & i_multiplicand[27];
wire w_pp_17_28 = i_multiplier[17] & i_multiplicand[28];
wire w_pp_17_29 = i_multiplier[17] & i_multiplicand[29];
wire w_pp_17_30 = i_multiplier[17] & i_multiplicand[30];
wire w_pp_17_31 = i_multiplier[17] & i_multiplicand[31];
wire w_pp_18_00 = i_multiplier[18] & i_multiplicand[ 0];
wire w_pp_18_01 = i_multiplier[18] & i_multiplicand[ 1];
wire w_pp_18_02 = i_multiplier[18] & i_multiplicand[ 2];
wire w_pp_18_03 = i_multiplier[18] & i_multiplicand[ 3];
wire w_pp_18_04 = i_multiplier[18] & i_multiplicand[ 4];
wire w_pp_18_05 = i_multiplier[18] & i_multiplicand[ 5];
wire w_pp_18_06 = i_multiplier[18] & i_multiplicand[ 6];
wire w_pp_18_07 = i_multiplier[18] & i_multiplicand[ 7];
wire w_pp_18_08 = i_multiplier[18] & i_multiplicand[ 8];
wire w_pp_18_09 = i_multiplier[18] & i_multiplicand[ 9];
wire w_pp_18_10 = i_multiplier[18] & i_multiplicand[10];
wire w_pp_18_11 = i_multiplier[18] & i_multiplicand[11];
wire w_pp_18_12 = i_multiplier[18] & i_multiplicand[12];
wire w_pp_18_13 = i_multiplier[18] & i_multiplicand[13];
wire w_pp_18_14 = i_multiplier[18] & i_multiplicand[14];
wire w_pp_18_15 = i_multiplier[18] & i_multiplicand[15];
wire w_pp_18_16 = i_multiplier[18] & i_multiplicand[16];
wire w_pp_18_17 = i_multiplier[18] & i_multiplicand[17];
wire w_pp_18_18 = i_multiplier[18] & i_multiplicand[18];
wire w_pp_18_19 = i_multiplier[18] & i_multiplicand[19];
wire w_pp_18_20 = i_multiplier[18] & i_multiplicand[20];
wire w_pp_18_21 = i_multiplier[18] & i_multiplicand[21];
wire w_pp_18_22 = i_multiplier[18] & i_multiplicand[22];
wire w_pp_18_23 = i_multiplier[18] & i_multiplicand[23];
wire w_pp_18_24 = i_multiplier[18] & i_multiplicand[24];
wire w_pp_18_25 = i_multiplier[18] & i_multiplicand[25];
wire w_pp_18_26 = i_multiplier[18] & i_multiplicand[26];
wire w_pp_18_27 = i_multiplier[18] & i_multiplicand[27];
wire w_pp_18_28 = i_multiplier[18] & i_multiplicand[28];
wire w_pp_18_29 = i_multiplier[18] & i_multiplicand[29];
wire w_pp_18_30 = i_multiplier[18] & i_multiplicand[30];
wire w_pp_18_31 = i_multiplier[18] & i_multiplicand[31];
wire w_pp_19_00 = i_multiplier[19] & i_multiplicand[ 0];
wire w_pp_19_01 = i_multiplier[19] & i_multiplicand[ 1];
wire w_pp_19_02 = i_multiplier[19] & i_multiplicand[ 2];
wire w_pp_19_03 = i_multiplier[19] & i_multiplicand[ 3];
wire w_pp_19_04 = i_multiplier[19] & i_multiplicand[ 4];
wire w_pp_19_05 = i_multiplier[19] & i_multiplicand[ 5];
wire w_pp_19_06 = i_multiplier[19] & i_multiplicand[ 6];
wire w_pp_19_07 = i_multiplier[19] & i_multiplicand[ 7];
wire w_pp_19_08 = i_multiplier[19] & i_multiplicand[ 8];
wire w_pp_19_09 = i_multiplier[19] & i_multiplicand[ 9];
wire w_pp_19_10 = i_multiplier[19] & i_multiplicand[10];
wire w_pp_19_11 = i_multiplier[19] & i_multiplicand[11];
wire w_pp_19_12 = i_multiplier[19] & i_multiplicand[12];
wire w_pp_19_13 = i_multiplier[19] & i_multiplicand[13];
wire w_pp_19_14 = i_multiplier[19] & i_multiplicand[14];
wire w_pp_19_15 = i_multiplier[19] & i_multiplicand[15];
wire w_pp_19_16 = i_multiplier[19] & i_multiplicand[16];
wire w_pp_19_17 = i_multiplier[19] & i_multiplicand[17];
wire w_pp_19_18 = i_multiplier[19] & i_multiplicand[18];
wire w_pp_19_19 = i_multiplier[19] & i_multiplicand[19];
wire w_pp_19_20 = i_multiplier[19] & i_multiplicand[20];
wire w_pp_19_21 = i_multiplier[19] & i_multiplicand[21];
wire w_pp_19_22 = i_multiplier[19] & i_multiplicand[22];
wire w_pp_19_23 = i_multiplier[19] & i_multiplicand[23];
wire w_pp_19_24 = i_multiplier[19] & i_multiplicand[24];
wire w_pp_19_25 = i_multiplier[19] & i_multiplicand[25];
wire w_pp_19_26 = i_multiplier[19] & i_multiplicand[26];
wire w_pp_19_27 = i_multiplier[19] & i_multiplicand[27];
wire w_pp_19_28 = i_multiplier[19] & i_multiplicand[28];
wire w_pp_19_29 = i_multiplier[19] & i_multiplicand[29];
wire w_pp_19_30 = i_multiplier[19] & i_multiplicand[30];
wire w_pp_19_31 = i_multiplier[19] & i_multiplicand[31];
wire w_pp_20_00 = i_multiplier[20] & i_multiplicand[ 0];
wire w_pp_20_01 = i_multiplier[20] & i_multiplicand[ 1];
wire w_pp_20_02 = i_multiplier[20] & i_multiplicand[ 2];
wire w_pp_20_03 = i_multiplier[20] & i_multiplicand[ 3];
wire w_pp_20_04 = i_multiplier[20] & i_multiplicand[ 4];
wire w_pp_20_05 = i_multiplier[20] & i_multiplicand[ 5];
wire w_pp_20_06 = i_multiplier[20] & i_multiplicand[ 6];
wire w_pp_20_07 = i_multiplier[20] & i_multiplicand[ 7];
wire w_pp_20_08 = i_multiplier[20] & i_multiplicand[ 8];
wire w_pp_20_09 = i_multiplier[20] & i_multiplicand[ 9];
wire w_pp_20_10 = i_multiplier[20] & i_multiplicand[10];
wire w_pp_20_11 = i_multiplier[20] & i_multiplicand[11];
wire w_pp_20_12 = i_multiplier[20] & i_multiplicand[12];
wire w_pp_20_13 = i_multiplier[20] & i_multiplicand[13];
wire w_pp_20_14 = i_multiplier[20] & i_multiplicand[14];
wire w_pp_20_15 = i_multiplier[20] & i_multiplicand[15];
wire w_pp_20_16 = i_multiplier[20] & i_multiplicand[16];
wire w_pp_20_17 = i_multiplier[20] & i_multiplicand[17];
wire w_pp_20_18 = i_multiplier[20] & i_multiplicand[18];
wire w_pp_20_19 = i_multiplier[20] & i_multiplicand[19];
wire w_pp_20_20 = i_multiplier[20] & i_multiplicand[20];
wire w_pp_20_21 = i_multiplier[20] & i_multiplicand[21];
wire w_pp_20_22 = i_multiplier[20] & i_multiplicand[22];
wire w_pp_20_23 = i_multiplier[20] & i_multiplicand[23];
wire w_pp_20_24 = i_multiplier[20] & i_multiplicand[24];
wire w_pp_20_25 = i_multiplier[20] & i_multiplicand[25];
wire w_pp_20_26 = i_multiplier[20] & i_multiplicand[26];
wire w_pp_20_27 = i_multiplier[20] & i_multiplicand[27];
wire w_pp_20_28 = i_multiplier[20] & i_multiplicand[28];
wire w_pp_20_29 = i_multiplier[20] & i_multiplicand[29];
wire w_pp_20_30 = i_multiplier[20] & i_multiplicand[30];
wire w_pp_20_31 = i_multiplier[20] & i_multiplicand[31];
wire w_pp_21_00 = i_multiplier[21] & i_multiplicand[ 0];
wire w_pp_21_01 = i_multiplier[21] & i_multiplicand[ 1];
wire w_pp_21_02 = i_multiplier[21] & i_multiplicand[ 2];
wire w_pp_21_03 = i_multiplier[21] & i_multiplicand[ 3];
wire w_pp_21_04 = i_multiplier[21] & i_multiplicand[ 4];
wire w_pp_21_05 = i_multiplier[21] & i_multiplicand[ 5];
wire w_pp_21_06 = i_multiplier[21] & i_multiplicand[ 6];
wire w_pp_21_07 = i_multiplier[21] & i_multiplicand[ 7];
wire w_pp_21_08 = i_multiplier[21] & i_multiplicand[ 8];
wire w_pp_21_09 = i_multiplier[21] & i_multiplicand[ 9];
wire w_pp_21_10 = i_multiplier[21] & i_multiplicand[10];
wire w_pp_21_11 = i_multiplier[21] & i_multiplicand[11];
wire w_pp_21_12 = i_multiplier[21] & i_multiplicand[12];
wire w_pp_21_13 = i_multiplier[21] & i_multiplicand[13];
wire w_pp_21_14 = i_multiplier[21] & i_multiplicand[14];
wire w_pp_21_15 = i_multiplier[21] & i_multiplicand[15];
wire w_pp_21_16 = i_multiplier[21] & i_multiplicand[16];
wire w_pp_21_17 = i_multiplier[21] & i_multiplicand[17];
wire w_pp_21_18 = i_multiplier[21] & i_multiplicand[18];
wire w_pp_21_19 = i_multiplier[21] & i_multiplicand[19];
wire w_pp_21_20 = i_multiplier[21] & i_multiplicand[20];
wire w_pp_21_21 = i_multiplier[21] & i_multiplicand[21];
wire w_pp_21_22 = i_multiplier[21] & i_multiplicand[22];
wire w_pp_21_23 = i_multiplier[21] & i_multiplicand[23];
wire w_pp_21_24 = i_multiplier[21] & i_multiplicand[24];
wire w_pp_21_25 = i_multiplier[21] & i_multiplicand[25];
wire w_pp_21_26 = i_multiplier[21] & i_multiplicand[26];
wire w_pp_21_27 = i_multiplier[21] & i_multiplicand[27];
wire w_pp_21_28 = i_multiplier[21] & i_multiplicand[28];
wire w_pp_21_29 = i_multiplier[21] & i_multiplicand[29];
wire w_pp_21_30 = i_multiplier[21] & i_multiplicand[30];
wire w_pp_21_31 = i_multiplier[21] & i_multiplicand[31];
wire w_pp_22_00 = i_multiplier[22] & i_multiplicand[ 0];
wire w_pp_22_01 = i_multiplier[22] & i_multiplicand[ 1];
wire w_pp_22_02 = i_multiplier[22] & i_multiplicand[ 2];
wire w_pp_22_03 = i_multiplier[22] & i_multiplicand[ 3];
wire w_pp_22_04 = i_multiplier[22] & i_multiplicand[ 4];
wire w_pp_22_05 = i_multiplier[22] & i_multiplicand[ 5];
wire w_pp_22_06 = i_multiplier[22] & i_multiplicand[ 6];
wire w_pp_22_07 = i_multiplier[22] & i_multiplicand[ 7];
wire w_pp_22_08 = i_multiplier[22] & i_multiplicand[ 8];
wire w_pp_22_09 = i_multiplier[22] & i_multiplicand[ 9];
wire w_pp_22_10 = i_multiplier[22] & i_multiplicand[10];
wire w_pp_22_11 = i_multiplier[22] & i_multiplicand[11];
wire w_pp_22_12 = i_multiplier[22] & i_multiplicand[12];
wire w_pp_22_13 = i_multiplier[22] & i_multiplicand[13];
wire w_pp_22_14 = i_multiplier[22] & i_multiplicand[14];
wire w_pp_22_15 = i_multiplier[22] & i_multiplicand[15];
wire w_pp_22_16 = i_multiplier[22] & i_multiplicand[16];
wire w_pp_22_17 = i_multiplier[22] & i_multiplicand[17];
wire w_pp_22_18 = i_multiplier[22] & i_multiplicand[18];
wire w_pp_22_19 = i_multiplier[22] & i_multiplicand[19];
wire w_pp_22_20 = i_multiplier[22] & i_multiplicand[20];
wire w_pp_22_21 = i_multiplier[22] & i_multiplicand[21];
wire w_pp_22_22 = i_multiplier[22] & i_multiplicand[22];
wire w_pp_22_23 = i_multiplier[22] & i_multiplicand[23];
wire w_pp_22_24 = i_multiplier[22] & i_multiplicand[24];
wire w_pp_22_25 = i_multiplier[22] & i_multiplicand[25];
wire w_pp_22_26 = i_multiplier[22] & i_multiplicand[26];
wire w_pp_22_27 = i_multiplier[22] & i_multiplicand[27];
wire w_pp_22_28 = i_multiplier[22] & i_multiplicand[28];
wire w_pp_22_29 = i_multiplier[22] & i_multiplicand[29];
wire w_pp_22_30 = i_multiplier[22] & i_multiplicand[30];
wire w_pp_22_31 = i_multiplier[22] & i_multiplicand[31];
wire w_pp_23_00 = i_multiplier[23] & i_multiplicand[ 0];
wire w_pp_23_01 = i_multiplier[23] & i_multiplicand[ 1];
wire w_pp_23_02 = i_multiplier[23] & i_multiplicand[ 2];
wire w_pp_23_03 = i_multiplier[23] & i_multiplicand[ 3];
wire w_pp_23_04 = i_multiplier[23] & i_multiplicand[ 4];
wire w_pp_23_05 = i_multiplier[23] & i_multiplicand[ 5];
wire w_pp_23_06 = i_multiplier[23] & i_multiplicand[ 6];
wire w_pp_23_07 = i_multiplier[23] & i_multiplicand[ 7];
wire w_pp_23_08 = i_multiplier[23] & i_multiplicand[ 8];
wire w_pp_23_09 = i_multiplier[23] & i_multiplicand[ 9];
wire w_pp_23_10 = i_multiplier[23] & i_multiplicand[10];
wire w_pp_23_11 = i_multiplier[23] & i_multiplicand[11];
wire w_pp_23_12 = i_multiplier[23] & i_multiplicand[12];
wire w_pp_23_13 = i_multiplier[23] & i_multiplicand[13];
wire w_pp_23_14 = i_multiplier[23] & i_multiplicand[14];
wire w_pp_23_15 = i_multiplier[23] & i_multiplicand[15];
wire w_pp_23_16 = i_multiplier[23] & i_multiplicand[16];
wire w_pp_23_17 = i_multiplier[23] & i_multiplicand[17];
wire w_pp_23_18 = i_multiplier[23] & i_multiplicand[18];
wire w_pp_23_19 = i_multiplier[23] & i_multiplicand[19];
wire w_pp_23_20 = i_multiplier[23] & i_multiplicand[20];
wire w_pp_23_21 = i_multiplier[23] & i_multiplicand[21];
wire w_pp_23_22 = i_multiplier[23] & i_multiplicand[22];
wire w_pp_23_23 = i_multiplier[23] & i_multiplicand[23];
wire w_pp_23_24 = i_multiplier[23] & i_multiplicand[24];
wire w_pp_23_25 = i_multiplier[23] & i_multiplicand[25];
wire w_pp_23_26 = i_multiplier[23] & i_multiplicand[26];
wire w_pp_23_27 = i_multiplier[23] & i_multiplicand[27];
wire w_pp_23_28 = i_multiplier[23] & i_multiplicand[28];
wire w_pp_23_29 = i_multiplier[23] & i_multiplicand[29];
wire w_pp_23_30 = i_multiplier[23] & i_multiplicand[30];
wire w_pp_23_31 = i_multiplier[23] & i_multiplicand[31];
wire w_pp_24_00 = i_multiplier[24] & i_multiplicand[ 0];
wire w_pp_24_01 = i_multiplier[24] & i_multiplicand[ 1];
wire w_pp_24_02 = i_multiplier[24] & i_multiplicand[ 2];
wire w_pp_24_03 = i_multiplier[24] & i_multiplicand[ 3];
wire w_pp_24_04 = i_multiplier[24] & i_multiplicand[ 4];
wire w_pp_24_05 = i_multiplier[24] & i_multiplicand[ 5];
wire w_pp_24_06 = i_multiplier[24] & i_multiplicand[ 6];
wire w_pp_24_07 = i_multiplier[24] & i_multiplicand[ 7];
wire w_pp_24_08 = i_multiplier[24] & i_multiplicand[ 8];
wire w_pp_24_09 = i_multiplier[24] & i_multiplicand[ 9];
wire w_pp_24_10 = i_multiplier[24] & i_multiplicand[10];
wire w_pp_24_11 = i_multiplier[24] & i_multiplicand[11];
wire w_pp_24_12 = i_multiplier[24] & i_multiplicand[12];
wire w_pp_24_13 = i_multiplier[24] & i_multiplicand[13];
wire w_pp_24_14 = i_multiplier[24] & i_multiplicand[14];
wire w_pp_24_15 = i_multiplier[24] & i_multiplicand[15];
wire w_pp_24_16 = i_multiplier[24] & i_multiplicand[16];
wire w_pp_24_17 = i_multiplier[24] & i_multiplicand[17];
wire w_pp_24_18 = i_multiplier[24] & i_multiplicand[18];
wire w_pp_24_19 = i_multiplier[24] & i_multiplicand[19];
wire w_pp_24_20 = i_multiplier[24] & i_multiplicand[20];
wire w_pp_24_21 = i_multiplier[24] & i_multiplicand[21];
wire w_pp_24_22 = i_multiplier[24] & i_multiplicand[22];
wire w_pp_24_23 = i_multiplier[24] & i_multiplicand[23];
wire w_pp_24_24 = i_multiplier[24] & i_multiplicand[24];
wire w_pp_24_25 = i_multiplier[24] & i_multiplicand[25];
wire w_pp_24_26 = i_multiplier[24] & i_multiplicand[26];
wire w_pp_24_27 = i_multiplier[24] & i_multiplicand[27];
wire w_pp_24_28 = i_multiplier[24] & i_multiplicand[28];
wire w_pp_24_29 = i_multiplier[24] & i_multiplicand[29];
wire w_pp_24_30 = i_multiplier[24] & i_multiplicand[30];
wire w_pp_24_31 = i_multiplier[24] & i_multiplicand[31];
wire w_pp_25_00 = i_multiplier[25] & i_multiplicand[ 0];
wire w_pp_25_01 = i_multiplier[25] & i_multiplicand[ 1];
wire w_pp_25_02 = i_multiplier[25] & i_multiplicand[ 2];
wire w_pp_25_03 = i_multiplier[25] & i_multiplicand[ 3];
wire w_pp_25_04 = i_multiplier[25] & i_multiplicand[ 4];
wire w_pp_25_05 = i_multiplier[25] & i_multiplicand[ 5];
wire w_pp_25_06 = i_multiplier[25] & i_multiplicand[ 6];
wire w_pp_25_07 = i_multiplier[25] & i_multiplicand[ 7];
wire w_pp_25_08 = i_multiplier[25] & i_multiplicand[ 8];
wire w_pp_25_09 = i_multiplier[25] & i_multiplicand[ 9];
wire w_pp_25_10 = i_multiplier[25] & i_multiplicand[10];
wire w_pp_25_11 = i_multiplier[25] & i_multiplicand[11];
wire w_pp_25_12 = i_multiplier[25] & i_multiplicand[12];
wire w_pp_25_13 = i_multiplier[25] & i_multiplicand[13];
wire w_pp_25_14 = i_multiplier[25] & i_multiplicand[14];
wire w_pp_25_15 = i_multiplier[25] & i_multiplicand[15];
wire w_pp_25_16 = i_multiplier[25] & i_multiplicand[16];
wire w_pp_25_17 = i_multiplier[25] & i_multiplicand[17];
wire w_pp_25_18 = i_multiplier[25] & i_multiplicand[18];
wire w_pp_25_19 = i_multiplier[25] & i_multiplicand[19];
wire w_pp_25_20 = i_multiplier[25] & i_multiplicand[20];
wire w_pp_25_21 = i_multiplier[25] & i_multiplicand[21];
wire w_pp_25_22 = i_multiplier[25] & i_multiplicand[22];
wire w_pp_25_23 = i_multiplier[25] & i_multiplicand[23];
wire w_pp_25_24 = i_multiplier[25] & i_multiplicand[24];
wire w_pp_25_25 = i_multiplier[25] & i_multiplicand[25];
wire w_pp_25_26 = i_multiplier[25] & i_multiplicand[26];
wire w_pp_25_27 = i_multiplier[25] & i_multiplicand[27];
wire w_pp_25_28 = i_multiplier[25] & i_multiplicand[28];
wire w_pp_25_29 = i_multiplier[25] & i_multiplicand[29];
wire w_pp_25_30 = i_multiplier[25] & i_multiplicand[30];
wire w_pp_25_31 = i_multiplier[25] & i_multiplicand[31];
wire w_pp_26_00 = i_multiplier[26] & i_multiplicand[ 0];
wire w_pp_26_01 = i_multiplier[26] & i_multiplicand[ 1];
wire w_pp_26_02 = i_multiplier[26] & i_multiplicand[ 2];
wire w_pp_26_03 = i_multiplier[26] & i_multiplicand[ 3];
wire w_pp_26_04 = i_multiplier[26] & i_multiplicand[ 4];
wire w_pp_26_05 = i_multiplier[26] & i_multiplicand[ 5];
wire w_pp_26_06 = i_multiplier[26] & i_multiplicand[ 6];
wire w_pp_26_07 = i_multiplier[26] & i_multiplicand[ 7];
wire w_pp_26_08 = i_multiplier[26] & i_multiplicand[ 8];
wire w_pp_26_09 = i_multiplier[26] & i_multiplicand[ 9];
wire w_pp_26_10 = i_multiplier[26] & i_multiplicand[10];
wire w_pp_26_11 = i_multiplier[26] & i_multiplicand[11];
wire w_pp_26_12 = i_multiplier[26] & i_multiplicand[12];
wire w_pp_26_13 = i_multiplier[26] & i_multiplicand[13];
wire w_pp_26_14 = i_multiplier[26] & i_multiplicand[14];
wire w_pp_26_15 = i_multiplier[26] & i_multiplicand[15];
wire w_pp_26_16 = i_multiplier[26] & i_multiplicand[16];
wire w_pp_26_17 = i_multiplier[26] & i_multiplicand[17];
wire w_pp_26_18 = i_multiplier[26] & i_multiplicand[18];
wire w_pp_26_19 = i_multiplier[26] & i_multiplicand[19];
wire w_pp_26_20 = i_multiplier[26] & i_multiplicand[20];
wire w_pp_26_21 = i_multiplier[26] & i_multiplicand[21];
wire w_pp_26_22 = i_multiplier[26] & i_multiplicand[22];
wire w_pp_26_23 = i_multiplier[26] & i_multiplicand[23];
wire w_pp_26_24 = i_multiplier[26] & i_multiplicand[24];
wire w_pp_26_25 = i_multiplier[26] & i_multiplicand[25];
wire w_pp_26_26 = i_multiplier[26] & i_multiplicand[26];
wire w_pp_26_27 = i_multiplier[26] & i_multiplicand[27];
wire w_pp_26_28 = i_multiplier[26] & i_multiplicand[28];
wire w_pp_26_29 = i_multiplier[26] & i_multiplicand[29];
wire w_pp_26_30 = i_multiplier[26] & i_multiplicand[30];
wire w_pp_26_31 = i_multiplier[26] & i_multiplicand[31];
wire w_pp_27_00 = i_multiplier[27] & i_multiplicand[ 0];
wire w_pp_27_01 = i_multiplier[27] & i_multiplicand[ 1];
wire w_pp_27_02 = i_multiplier[27] & i_multiplicand[ 2];
wire w_pp_27_03 = i_multiplier[27] & i_multiplicand[ 3];
wire w_pp_27_04 = i_multiplier[27] & i_multiplicand[ 4];
wire w_pp_27_05 = i_multiplier[27] & i_multiplicand[ 5];
wire w_pp_27_06 = i_multiplier[27] & i_multiplicand[ 6];
wire w_pp_27_07 = i_multiplier[27] & i_multiplicand[ 7];
wire w_pp_27_08 = i_multiplier[27] & i_multiplicand[ 8];
wire w_pp_27_09 = i_multiplier[27] & i_multiplicand[ 9];
wire w_pp_27_10 = i_multiplier[27] & i_multiplicand[10];
wire w_pp_27_11 = i_multiplier[27] & i_multiplicand[11];
wire w_pp_27_12 = i_multiplier[27] & i_multiplicand[12];
wire w_pp_27_13 = i_multiplier[27] & i_multiplicand[13];
wire w_pp_27_14 = i_multiplier[27] & i_multiplicand[14];
wire w_pp_27_15 = i_multiplier[27] & i_multiplicand[15];
wire w_pp_27_16 = i_multiplier[27] & i_multiplicand[16];
wire w_pp_27_17 = i_multiplier[27] & i_multiplicand[17];
wire w_pp_27_18 = i_multiplier[27] & i_multiplicand[18];
wire w_pp_27_19 = i_multiplier[27] & i_multiplicand[19];
wire w_pp_27_20 = i_multiplier[27] & i_multiplicand[20];
wire w_pp_27_21 = i_multiplier[27] & i_multiplicand[21];
wire w_pp_27_22 = i_multiplier[27] & i_multiplicand[22];
wire w_pp_27_23 = i_multiplier[27] & i_multiplicand[23];
wire w_pp_27_24 = i_multiplier[27] & i_multiplicand[24];
wire w_pp_27_25 = i_multiplier[27] & i_multiplicand[25];
wire w_pp_27_26 = i_multiplier[27] & i_multiplicand[26];
wire w_pp_27_27 = i_multiplier[27] & i_multiplicand[27];
wire w_pp_27_28 = i_multiplier[27] & i_multiplicand[28];
wire w_pp_27_29 = i_multiplier[27] & i_multiplicand[29];
wire w_pp_27_30 = i_multiplier[27] & i_multiplicand[30];
wire w_pp_27_31 = i_multiplier[27] & i_multiplicand[31];
wire w_pp_28_00 = i_multiplier[28] & i_multiplicand[ 0];
wire w_pp_28_01 = i_multiplier[28] & i_multiplicand[ 1];
wire w_pp_28_02 = i_multiplier[28] & i_multiplicand[ 2];
wire w_pp_28_03 = i_multiplier[28] & i_multiplicand[ 3];
wire w_pp_28_04 = i_multiplier[28] & i_multiplicand[ 4];
wire w_pp_28_05 = i_multiplier[28] & i_multiplicand[ 5];
wire w_pp_28_06 = i_multiplier[28] & i_multiplicand[ 6];
wire w_pp_28_07 = i_multiplier[28] & i_multiplicand[ 7];
wire w_pp_28_08 = i_multiplier[28] & i_multiplicand[ 8];
wire w_pp_28_09 = i_multiplier[28] & i_multiplicand[ 9];
wire w_pp_28_10 = i_multiplier[28] & i_multiplicand[10];
wire w_pp_28_11 = i_multiplier[28] & i_multiplicand[11];
wire w_pp_28_12 = i_multiplier[28] & i_multiplicand[12];
wire w_pp_28_13 = i_multiplier[28] & i_multiplicand[13];
wire w_pp_28_14 = i_multiplier[28] & i_multiplicand[14];
wire w_pp_28_15 = i_multiplier[28] & i_multiplicand[15];
wire w_pp_28_16 = i_multiplier[28] & i_multiplicand[16];
wire w_pp_28_17 = i_multiplier[28] & i_multiplicand[17];
wire w_pp_28_18 = i_multiplier[28] & i_multiplicand[18];
wire w_pp_28_19 = i_multiplier[28] & i_multiplicand[19];
wire w_pp_28_20 = i_multiplier[28] & i_multiplicand[20];
wire w_pp_28_21 = i_multiplier[28] & i_multiplicand[21];
wire w_pp_28_22 = i_multiplier[28] & i_multiplicand[22];
wire w_pp_28_23 = i_multiplier[28] & i_multiplicand[23];
wire w_pp_28_24 = i_multiplier[28] & i_multiplicand[24];
wire w_pp_28_25 = i_multiplier[28] & i_multiplicand[25];
wire w_pp_28_26 = i_multiplier[28] & i_multiplicand[26];
wire w_pp_28_27 = i_multiplier[28] & i_multiplicand[27];
wire w_pp_28_28 = i_multiplier[28] & i_multiplicand[28];
wire w_pp_28_29 = i_multiplier[28] & i_multiplicand[29];
wire w_pp_28_30 = i_multiplier[28] & i_multiplicand[30];
wire w_pp_28_31 = i_multiplier[28] & i_multiplicand[31];
wire w_pp_29_00 = i_multiplier[29] & i_multiplicand[ 0];
wire w_pp_29_01 = i_multiplier[29] & i_multiplicand[ 1];
wire w_pp_29_02 = i_multiplier[29] & i_multiplicand[ 2];
wire w_pp_29_03 = i_multiplier[29] & i_multiplicand[ 3];
wire w_pp_29_04 = i_multiplier[29] & i_multiplicand[ 4];
wire w_pp_29_05 = i_multiplier[29] & i_multiplicand[ 5];
wire w_pp_29_06 = i_multiplier[29] & i_multiplicand[ 6];
wire w_pp_29_07 = i_multiplier[29] & i_multiplicand[ 7];
wire w_pp_29_08 = i_multiplier[29] & i_multiplicand[ 8];
wire w_pp_29_09 = i_multiplier[29] & i_multiplicand[ 9];
wire w_pp_29_10 = i_multiplier[29] & i_multiplicand[10];
wire w_pp_29_11 = i_multiplier[29] & i_multiplicand[11];
wire w_pp_29_12 = i_multiplier[29] & i_multiplicand[12];
wire w_pp_29_13 = i_multiplier[29] & i_multiplicand[13];
wire w_pp_29_14 = i_multiplier[29] & i_multiplicand[14];
wire w_pp_29_15 = i_multiplier[29] & i_multiplicand[15];
wire w_pp_29_16 = i_multiplier[29] & i_multiplicand[16];
wire w_pp_29_17 = i_multiplier[29] & i_multiplicand[17];
wire w_pp_29_18 = i_multiplier[29] & i_multiplicand[18];
wire w_pp_29_19 = i_multiplier[29] & i_multiplicand[19];
wire w_pp_29_20 = i_multiplier[29] & i_multiplicand[20];
wire w_pp_29_21 = i_multiplier[29] & i_multiplicand[21];
wire w_pp_29_22 = i_multiplier[29] & i_multiplicand[22];
wire w_pp_29_23 = i_multiplier[29] & i_multiplicand[23];
wire w_pp_29_24 = i_multiplier[29] & i_multiplicand[24];
wire w_pp_29_25 = i_multiplier[29] & i_multiplicand[25];
wire w_pp_29_26 = i_multiplier[29] & i_multiplicand[26];
wire w_pp_29_27 = i_multiplier[29] & i_multiplicand[27];
wire w_pp_29_28 = i_multiplier[29] & i_multiplicand[28];
wire w_pp_29_29 = i_multiplier[29] & i_multiplicand[29];
wire w_pp_29_30 = i_multiplier[29] & i_multiplicand[30];
wire w_pp_29_31 = i_multiplier[29] & i_multiplicand[31];
wire w_pp_30_00 = i_multiplier[30] & i_multiplicand[ 0];
wire w_pp_30_01 = i_multiplier[30] & i_multiplicand[ 1];
wire w_pp_30_02 = i_multiplier[30] & i_multiplicand[ 2];
wire w_pp_30_03 = i_multiplier[30] & i_multiplicand[ 3];
wire w_pp_30_04 = i_multiplier[30] & i_multiplicand[ 4];
wire w_pp_30_05 = i_multiplier[30] & i_multiplicand[ 5];
wire w_pp_30_06 = i_multiplier[30] & i_multiplicand[ 6];
wire w_pp_30_07 = i_multiplier[30] & i_multiplicand[ 7];
wire w_pp_30_08 = i_multiplier[30] & i_multiplicand[ 8];
wire w_pp_30_09 = i_multiplier[30] & i_multiplicand[ 9];
wire w_pp_30_10 = i_multiplier[30] & i_multiplicand[10];
wire w_pp_30_11 = i_multiplier[30] & i_multiplicand[11];
wire w_pp_30_12 = i_multiplier[30] & i_multiplicand[12];
wire w_pp_30_13 = i_multiplier[30] & i_multiplicand[13];
wire w_pp_30_14 = i_multiplier[30] & i_multiplicand[14];
wire w_pp_30_15 = i_multiplier[30] & i_multiplicand[15];
wire w_pp_30_16 = i_multiplier[30] & i_multiplicand[16];
wire w_pp_30_17 = i_multiplier[30] & i_multiplicand[17];
wire w_pp_30_18 = i_multiplier[30] & i_multiplicand[18];
wire w_pp_30_19 = i_multiplier[30] & i_multiplicand[19];
wire w_pp_30_20 = i_multiplier[30] & i_multiplicand[20];
wire w_pp_30_21 = i_multiplier[30] & i_multiplicand[21];
wire w_pp_30_22 = i_multiplier[30] & i_multiplicand[22];
wire w_pp_30_23 = i_multiplier[30] & i_multiplicand[23];
wire w_pp_30_24 = i_multiplier[30] & i_multiplicand[24];
wire w_pp_30_25 = i_multiplier[30] & i_multiplicand[25];
wire w_pp_30_26 = i_multiplier[30] & i_multiplicand[26];
wire w_pp_30_27 = i_multiplier[30] & i_multiplicand[27];
wire w_pp_30_28 = i_multiplier[30] & i_multiplicand[28];
wire w_pp_30_29 = i_multiplier[30] & i_multiplicand[29];
wire w_pp_30_30 = i_multiplier[30] & i_multiplicand[30];
wire w_pp_30_31 = i_multiplier[30] & i_multiplicand[31];
wire w_pp_31_00 = i_multiplier[31] & i_multiplicand[ 0];
wire w_pp_31_01 = i_multiplier[31] & i_multiplicand[ 1];
wire w_pp_31_02 = i_multiplier[31] & i_multiplicand[ 2];
wire w_pp_31_03 = i_multiplier[31] & i_multiplicand[ 3];
wire w_pp_31_04 = i_multiplier[31] & i_multiplicand[ 4];
wire w_pp_31_05 = i_multiplier[31] & i_multiplicand[ 5];
wire w_pp_31_06 = i_multiplier[31] & i_multiplicand[ 6];
wire w_pp_31_07 = i_multiplier[31] & i_multiplicand[ 7];
wire w_pp_31_08 = i_multiplier[31] & i_multiplicand[ 8];
wire w_pp_31_09 = i_multiplier[31] & i_multiplicand[ 9];
wire w_pp_31_10 = i_multiplier[31] & i_multiplicand[10];
wire w_pp_31_11 = i_multiplier[31] & i_multiplicand[11];
wire w_pp_31_12 = i_multiplier[31] & i_multiplicand[12];
wire w_pp_31_13 = i_multiplier[31] & i_multiplicand[13];
wire w_pp_31_14 = i_multiplier[31] & i_multiplicand[14];
wire w_pp_31_15 = i_multiplier[31] & i_multiplicand[15];
wire w_pp_31_16 = i_multiplier[31] & i_multiplicand[16];
wire w_pp_31_17 = i_multiplier[31] & i_multiplicand[17];
wire w_pp_31_18 = i_multiplier[31] & i_multiplicand[18];
wire w_pp_31_19 = i_multiplier[31] & i_multiplicand[19];
wire w_pp_31_20 = i_multiplier[31] & i_multiplicand[20];
wire w_pp_31_21 = i_multiplier[31] & i_multiplicand[21];
wire w_pp_31_22 = i_multiplier[31] & i_multiplicand[22];
wire w_pp_31_23 = i_multiplier[31] & i_multiplicand[23];
wire w_pp_31_24 = i_multiplier[31] & i_multiplicand[24];
wire w_pp_31_25 = i_multiplier[31] & i_multiplicand[25];
wire w_pp_31_26 = i_multiplier[31] & i_multiplicand[26];
wire w_pp_31_27 = i_multiplier[31] & i_multiplicand[27];
wire w_pp_31_28 = i_multiplier[31] & i_multiplicand[28];
wire w_pp_31_29 = i_multiplier[31] & i_multiplicand[29];
wire w_pp_31_30 = i_multiplier[31] & i_multiplicand[30];
wire w_pp_31_31 = i_multiplier[31] & i_multiplicand[31];

// Stage: 0, Max Height: 24
wire w_sum_0, w_carry_0;
math_adder_half HA_0(.i_a(w_pp_00_24), .i_b(w_pp_01_23), .ow_sum(w_sum_0), .ow_carry(w_carry_0));
wire w_sum_1, w_carry_1;
math_adder_carry_save CSA_1(.i_a(w_pp_00_25), .i_b(w_pp_01_24), .i_c(w_pp_02_23), .ow_sum(w_sum_1), .ow_carry(w_carry_1));
wire w_sum_2, w_carry_2;
math_adder_half HA_2(.i_a(w_pp_03_22), .i_b(w_pp_04_21), .ow_sum(w_sum_2), .ow_carry(w_carry_2));
wire w_sum_3, w_carry_3;
math_adder_carry_save CSA_3(.i_a(w_pp_00_26), .i_b(w_pp_01_25), .i_c(w_pp_02_24), .ow_sum(w_sum_3), .ow_carry(w_carry_3));
wire w_sum_4, w_carry_4;
math_adder_carry_save CSA_4(.i_a(w_pp_03_23), .i_b(w_pp_04_22), .i_c(w_pp_05_21), .ow_sum(w_sum_4), .ow_carry(w_carry_4));
wire w_sum_5, w_carry_5;
math_adder_half HA_5(.i_a(w_pp_06_20), .i_b(w_pp_07_19), .ow_sum(w_sum_5), .ow_carry(w_carry_5));
wire w_sum_6, w_carry_6;
math_adder_carry_save CSA_6(.i_a(w_pp_00_27), .i_b(w_pp_01_26), .i_c(w_pp_02_25), .ow_sum(w_sum_6), .ow_carry(w_carry_6));
wire w_sum_7, w_carry_7;
math_adder_carry_save CSA_7(.i_a(w_pp_03_24), .i_b(w_pp_04_23), .i_c(w_pp_05_22), .ow_sum(w_sum_7), .ow_carry(w_carry_7));
wire w_sum_8, w_carry_8;
math_adder_carry_save CSA_8(.i_a(w_pp_06_21), .i_b(w_pp_07_20), .i_c(w_pp_08_19), .ow_sum(w_sum_8), .ow_carry(w_carry_8));
wire w_sum_9, w_carry_9;
math_adder_half HA_9(.i_a(w_pp_09_18), .i_b(w_pp_10_17), .ow_sum(w_sum_9), .ow_carry(w_carry_9));
wire w_sum_10, w_carry_10;
math_adder_carry_save CSA_10(.i_a(w_pp_00_28), .i_b(w_pp_01_27), .i_c(w_pp_02_26), .ow_sum(w_sum_10), .ow_carry(w_carry_10));
wire w_sum_11, w_carry_11;
math_adder_carry_save CSA_11(.i_a(w_pp_03_25), .i_b(w_pp_04_24), .i_c(w_pp_05_23), .ow_sum(w_sum_11), .ow_carry(w_carry_11));
wire w_sum_12, w_carry_12;
math_adder_carry_save CSA_12(.i_a(w_pp_06_22), .i_b(w_pp_07_21), .i_c(w_pp_08_20), .ow_sum(w_sum_12), .ow_carry(w_carry_12));
wire w_sum_13, w_carry_13;
math_adder_carry_save CSA_13(.i_a(w_pp_09_19), .i_b(w_pp_10_18), .i_c(w_pp_11_17), .ow_sum(w_sum_13), .ow_carry(w_carry_13));
wire w_sum_14, w_carry_14;
math_adder_half HA_14(.i_a(w_pp_12_16), .i_b(w_pp_13_15), .ow_sum(w_sum_14), .ow_carry(w_carry_14));
wire w_sum_15, w_carry_15;
math_adder_carry_save CSA_15(.i_a(w_pp_00_29), .i_b(w_pp_01_28), .i_c(w_pp_02_27), .ow_sum(w_sum_15), .ow_carry(w_carry_15));
wire w_sum_16, w_carry_16;
math_adder_carry_save CSA_16(.i_a(w_pp_03_26), .i_b(w_pp_04_25), .i_c(w_pp_05_24), .ow_sum(w_sum_16), .ow_carry(w_carry_16));
wire w_sum_17, w_carry_17;
math_adder_carry_save CSA_17(.i_a(w_pp_06_23), .i_b(w_pp_07_22), .i_c(w_pp_08_21), .ow_sum(w_sum_17), .ow_carry(w_carry_17));
wire w_sum_18, w_carry_18;
math_adder_carry_save CSA_18(.i_a(w_pp_09_20), .i_b(w_pp_10_19), .i_c(w_pp_11_18), .ow_sum(w_sum_18), .ow_carry(w_carry_18));
wire w_sum_19, w_carry_19;
math_adder_carry_save CSA_19(.i_a(w_pp_12_17), .i_b(w_pp_13_16), .i_c(w_pp_14_15), .ow_sum(w_sum_19), .ow_carry(w_carry_19));
wire w_sum_20, w_carry_20;
math_adder_half HA_20(.i_a(w_pp_15_14), .i_b(w_pp_16_13), .ow_sum(w_sum_20), .ow_carry(w_carry_20));
wire w_sum_21, w_carry_21;
math_adder_carry_save CSA_21(.i_a(w_pp_00_30), .i_b(w_pp_01_29), .i_c(w_pp_02_28), .ow_sum(w_sum_21), .ow_carry(w_carry_21));
wire w_sum_22, w_carry_22;
math_adder_carry_save CSA_22(.i_a(w_pp_03_27), .i_b(w_pp_04_26), .i_c(w_pp_05_25), .ow_sum(w_sum_22), .ow_carry(w_carry_22));
wire w_sum_23, w_carry_23;
math_adder_carry_save CSA_23(.i_a(w_pp_06_24), .i_b(w_pp_07_23), .i_c(w_pp_08_22), .ow_sum(w_sum_23), .ow_carry(w_carry_23));
wire w_sum_24, w_carry_24;
math_adder_carry_save CSA_24(.i_a(w_pp_09_21), .i_b(w_pp_10_20), .i_c(w_pp_11_19), .ow_sum(w_sum_24), .ow_carry(w_carry_24));
wire w_sum_25, w_carry_25;
math_adder_carry_save CSA_25(.i_a(w_pp_12_18), .i_b(w_pp_13_17), .i_c(w_pp_14_16), .ow_sum(w_sum_25), .ow_carry(w_carry_25));
wire w_sum_26, w_carry_26;
math_adder_carry_save CSA_26(.i_a(w_pp_15_15), .i_b(w_pp_16_14), .i_c(w_pp_17_13), .ow_sum(w_sum_26), .ow_carry(w_carry_26));
wire w_sum_27, w_carry_27;
math_adder_half HA_27(.i_a(w_pp_18_12), .i_b(w_pp_19_11), .ow_sum(w_sum_27), .ow_carry(w_carry_27));
wire w_sum_28, w_carry_28;
math_adder_carry_save CSA_28(.i_a(w_pp_00_31), .i_b(w_pp_01_30), .i_c(w_pp_02_29), .ow_sum(w_sum_28), .ow_carry(w_carry_28));
wire w_sum_29, w_carry_29;
math_adder_carry_save CSA_29(.i_a(w_pp_03_28), .i_b(w_pp_04_27), .i_c(w_pp_05_26), .ow_sum(w_sum_29), .ow_carry(w_carry_29));
wire w_sum_30, w_carry_30;
math_adder_carry_save CSA_30(.i_a(w_pp_06_25), .i_b(w_pp_07_24), .i_c(w_pp_08_23), .ow_sum(w_sum_30), .ow_carry(w_carry_30));
wire w_sum_31, w_carry_31;
math_adder_carry_save CSA_31(.i_a(w_pp_09_22), .i_b(w_pp_10_21), .i_c(w_pp_11_20), .ow_sum(w_sum_31), .ow_carry(w_carry_31));
wire w_sum_32, w_carry_32;
math_adder_carry_save CSA_32(.i_a(w_pp_12_19), .i_b(w_pp_13_18), .i_c(w_pp_14_17), .ow_sum(w_sum_32), .ow_carry(w_carry_32));
wire w_sum_33, w_carry_33;
math_adder_carry_save CSA_33(.i_a(w_pp_15_16), .i_b(w_pp_16_15), .i_c(w_pp_17_14), .ow_sum(w_sum_33), .ow_carry(w_carry_33));
wire w_sum_34, w_carry_34;
math_adder_carry_save CSA_34(.i_a(w_pp_18_13), .i_b(w_pp_19_12), .i_c(w_pp_20_11), .ow_sum(w_sum_34), .ow_carry(w_carry_34));
wire w_sum_35, w_carry_35;
math_adder_half HA_35(.i_a(w_pp_21_10), .i_b(w_pp_22_09), .ow_sum(w_sum_35), .ow_carry(w_carry_35));
wire w_sum_36, w_carry_36;
math_adder_carry_save CSA_36(.i_a(w_pp_01_31), .i_b(w_pp_02_30), .i_c(w_pp_03_29), .ow_sum(w_sum_36), .ow_carry(w_carry_36));
wire w_sum_37, w_carry_37;
math_adder_carry_save CSA_37(.i_a(w_pp_04_28), .i_b(w_pp_05_27), .i_c(w_pp_06_26), .ow_sum(w_sum_37), .ow_carry(w_carry_37));
wire w_sum_38, w_carry_38;
math_adder_carry_save CSA_38(.i_a(w_pp_07_25), .i_b(w_pp_08_24), .i_c(w_pp_09_23), .ow_sum(w_sum_38), .ow_carry(w_carry_38));
wire w_sum_39, w_carry_39;
math_adder_carry_save CSA_39(.i_a(w_pp_10_22), .i_b(w_pp_11_21), .i_c(w_pp_12_20), .ow_sum(w_sum_39), .ow_carry(w_carry_39));
wire w_sum_40, w_carry_40;
math_adder_carry_save CSA_40(.i_a(w_pp_13_19), .i_b(w_pp_14_18), .i_c(w_pp_15_17), .ow_sum(w_sum_40), .ow_carry(w_carry_40));
wire w_sum_41, w_carry_41;
math_adder_carry_save CSA_41(.i_a(w_pp_16_16), .i_b(w_pp_17_15), .i_c(w_pp_18_14), .ow_sum(w_sum_41), .ow_carry(w_carry_41));
wire w_sum_42, w_carry_42;
math_adder_carry_save CSA_42(.i_a(w_pp_19_13), .i_b(w_pp_20_12), .i_c(w_pp_21_11), .ow_sum(w_sum_42), .ow_carry(w_carry_42));
wire w_sum_43, w_carry_43;
math_adder_half HA_43(.i_a(w_pp_22_10), .i_b(w_pp_23_09), .ow_sum(w_sum_43), .ow_carry(w_carry_43));
wire w_sum_44, w_carry_44;
math_adder_carry_save CSA_44(.i_a(w_pp_02_31), .i_b(w_pp_03_30), .i_c(w_pp_04_29), .ow_sum(w_sum_44), .ow_carry(w_carry_44));
wire w_sum_45, w_carry_45;
math_adder_carry_save CSA_45(.i_a(w_pp_05_28), .i_b(w_pp_06_27), .i_c(w_pp_07_26), .ow_sum(w_sum_45), .ow_carry(w_carry_45));
wire w_sum_46, w_carry_46;
math_adder_carry_save CSA_46(.i_a(w_pp_08_25), .i_b(w_pp_09_24), .i_c(w_pp_10_23), .ow_sum(w_sum_46), .ow_carry(w_carry_46));
wire w_sum_47, w_carry_47;
math_adder_carry_save CSA_47(.i_a(w_pp_11_22), .i_b(w_pp_12_21), .i_c(w_pp_13_20), .ow_sum(w_sum_47), .ow_carry(w_carry_47));
wire w_sum_48, w_carry_48;
math_adder_carry_save CSA_48(.i_a(w_pp_14_19), .i_b(w_pp_15_18), .i_c(w_pp_16_17), .ow_sum(w_sum_48), .ow_carry(w_carry_48));
wire w_sum_49, w_carry_49;
math_adder_carry_save CSA_49(.i_a(w_pp_17_16), .i_b(w_pp_18_15), .i_c(w_pp_19_14), .ow_sum(w_sum_49), .ow_carry(w_carry_49));
wire w_sum_50, w_carry_50;
math_adder_carry_save CSA_50(.i_a(w_pp_20_13), .i_b(w_pp_21_12), .i_c(w_pp_22_11), .ow_sum(w_sum_50), .ow_carry(w_carry_50));
wire w_sum_51, w_carry_51;
math_adder_carry_save CSA_51(.i_a(w_pp_03_31), .i_b(w_pp_04_30), .i_c(w_pp_05_29), .ow_sum(w_sum_51), .ow_carry(w_carry_51));
wire w_sum_52, w_carry_52;
math_adder_carry_save CSA_52(.i_a(w_pp_06_28), .i_b(w_pp_07_27), .i_c(w_pp_08_26), .ow_sum(w_sum_52), .ow_carry(w_carry_52));
wire w_sum_53, w_carry_53;
math_adder_carry_save CSA_53(.i_a(w_pp_09_25), .i_b(w_pp_10_24), .i_c(w_pp_11_23), .ow_sum(w_sum_53), .ow_carry(w_carry_53));
wire w_sum_54, w_carry_54;
math_adder_carry_save CSA_54(.i_a(w_pp_12_22), .i_b(w_pp_13_21), .i_c(w_pp_14_20), .ow_sum(w_sum_54), .ow_carry(w_carry_54));
wire w_sum_55, w_carry_55;
math_adder_carry_save CSA_55(.i_a(w_pp_15_19), .i_b(w_pp_16_18), .i_c(w_pp_17_17), .ow_sum(w_sum_55), .ow_carry(w_carry_55));
wire w_sum_56, w_carry_56;
math_adder_carry_save CSA_56(.i_a(w_pp_18_16), .i_b(w_pp_19_15), .i_c(w_pp_20_14), .ow_sum(w_sum_56), .ow_carry(w_carry_56));
wire w_sum_57, w_carry_57;
math_adder_carry_save CSA_57(.i_a(w_pp_04_31), .i_b(w_pp_05_30), .i_c(w_pp_06_29), .ow_sum(w_sum_57), .ow_carry(w_carry_57));
wire w_sum_58, w_carry_58;
math_adder_carry_save CSA_58(.i_a(w_pp_07_28), .i_b(w_pp_08_27), .i_c(w_pp_09_26), .ow_sum(w_sum_58), .ow_carry(w_carry_58));
wire w_sum_59, w_carry_59;
math_adder_carry_save CSA_59(.i_a(w_pp_10_25), .i_b(w_pp_11_24), .i_c(w_pp_12_23), .ow_sum(w_sum_59), .ow_carry(w_carry_59));
wire w_sum_60, w_carry_60;
math_adder_carry_save CSA_60(.i_a(w_pp_13_22), .i_b(w_pp_14_21), .i_c(w_pp_15_20), .ow_sum(w_sum_60), .ow_carry(w_carry_60));
wire w_sum_61, w_carry_61;
math_adder_carry_save CSA_61(.i_a(w_pp_16_19), .i_b(w_pp_17_18), .i_c(w_pp_18_17), .ow_sum(w_sum_61), .ow_carry(w_carry_61));
wire w_sum_62, w_carry_62;
math_adder_carry_save CSA_62(.i_a(w_pp_05_31), .i_b(w_pp_06_30), .i_c(w_pp_07_29), .ow_sum(w_sum_62), .ow_carry(w_carry_62));
wire w_sum_63, w_carry_63;
math_adder_carry_save CSA_63(.i_a(w_pp_08_28), .i_b(w_pp_09_27), .i_c(w_pp_10_26), .ow_sum(w_sum_63), .ow_carry(w_carry_63));
wire w_sum_64, w_carry_64;
math_adder_carry_save CSA_64(.i_a(w_pp_11_25), .i_b(w_pp_12_24), .i_c(w_pp_13_23), .ow_sum(w_sum_64), .ow_carry(w_carry_64));
wire w_sum_65, w_carry_65;
math_adder_carry_save CSA_65(.i_a(w_pp_14_22), .i_b(w_pp_15_21), .i_c(w_pp_16_20), .ow_sum(w_sum_65), .ow_carry(w_carry_65));
wire w_sum_66, w_carry_66;
math_adder_carry_save CSA_66(.i_a(w_pp_06_31), .i_b(w_pp_07_30), .i_c(w_pp_08_29), .ow_sum(w_sum_66), .ow_carry(w_carry_66));
wire w_sum_67, w_carry_67;
math_adder_carry_save CSA_67(.i_a(w_pp_09_28), .i_b(w_pp_10_27), .i_c(w_pp_11_26), .ow_sum(w_sum_67), .ow_carry(w_carry_67));
wire w_sum_68, w_carry_68;
math_adder_carry_save CSA_68(.i_a(w_pp_12_25), .i_b(w_pp_13_24), .i_c(w_pp_14_23), .ow_sum(w_sum_68), .ow_carry(w_carry_68));
wire w_sum_69, w_carry_69;
math_adder_carry_save CSA_69(.i_a(w_pp_07_31), .i_b(w_pp_08_30), .i_c(w_pp_09_29), .ow_sum(w_sum_69), .ow_carry(w_carry_69));
wire w_sum_70, w_carry_70;
math_adder_carry_save CSA_70(.i_a(w_pp_10_28), .i_b(w_pp_11_27), .i_c(w_pp_12_26), .ow_sum(w_sum_70), .ow_carry(w_carry_70));
wire w_sum_71, w_carry_71;
math_adder_carry_save CSA_71(.i_a(w_pp_08_31), .i_b(w_pp_09_30), .i_c(w_pp_10_29), .ow_sum(w_sum_71), .ow_carry(w_carry_71));
// Stage: 1, Max Height: 16
wire w_sum_72, w_carry_72;
math_adder_half HA_72(.i_a(w_pp_00_16), .i_b(w_pp_01_15), .ow_sum(w_sum_72), .ow_carry(w_carry_72));
wire w_sum_73, w_carry_73;
math_adder_carry_save CSA_73(.i_a(w_pp_00_17), .i_b(w_pp_01_16), .i_c(w_pp_02_15), .ow_sum(w_sum_73), .ow_carry(w_carry_73));
wire w_sum_74, w_carry_74;
math_adder_half HA_74(.i_a(w_pp_03_14), .i_b(w_pp_04_13), .ow_sum(w_sum_74), .ow_carry(w_carry_74));
wire w_sum_75, w_carry_75;
math_adder_carry_save CSA_75(.i_a(w_pp_00_18), .i_b(w_pp_01_17), .i_c(w_pp_02_16), .ow_sum(w_sum_75), .ow_carry(w_carry_75));
wire w_sum_76, w_carry_76;
math_adder_carry_save CSA_76(.i_a(w_pp_03_15), .i_b(w_pp_04_14), .i_c(w_pp_05_13), .ow_sum(w_sum_76), .ow_carry(w_carry_76));
wire w_sum_77, w_carry_77;
math_adder_half HA_77(.i_a(w_pp_06_12), .i_b(w_pp_07_11), .ow_sum(w_sum_77), .ow_carry(w_carry_77));
wire w_sum_78, w_carry_78;
math_adder_carry_save CSA_78(.i_a(w_pp_00_19), .i_b(w_pp_01_18), .i_c(w_pp_02_17), .ow_sum(w_sum_78), .ow_carry(w_carry_78));
wire w_sum_79, w_carry_79;
math_adder_carry_save CSA_79(.i_a(w_pp_03_16), .i_b(w_pp_04_15), .i_c(w_pp_05_14), .ow_sum(w_sum_79), .ow_carry(w_carry_79));
wire w_sum_80, w_carry_80;
math_adder_carry_save CSA_80(.i_a(w_pp_06_13), .i_b(w_pp_07_12), .i_c(w_pp_08_11), .ow_sum(w_sum_80), .ow_carry(w_carry_80));
wire w_sum_81, w_carry_81;
math_adder_half HA_81(.i_a(w_pp_09_10), .i_b(w_pp_10_09), .ow_sum(w_sum_81), .ow_carry(w_carry_81));
wire w_sum_82, w_carry_82;
math_adder_carry_save CSA_82(.i_a(w_pp_00_20), .i_b(w_pp_01_19), .i_c(w_pp_02_18), .ow_sum(w_sum_82), .ow_carry(w_carry_82));
wire w_sum_83, w_carry_83;
math_adder_carry_save CSA_83(.i_a(w_pp_03_17), .i_b(w_pp_04_16), .i_c(w_pp_05_15), .ow_sum(w_sum_83), .ow_carry(w_carry_83));
wire w_sum_84, w_carry_84;
math_adder_carry_save CSA_84(.i_a(w_pp_06_14), .i_b(w_pp_07_13), .i_c(w_pp_08_12), .ow_sum(w_sum_84), .ow_carry(w_carry_84));
wire w_sum_85, w_carry_85;
math_adder_carry_save CSA_85(.i_a(w_pp_09_11), .i_b(w_pp_10_10), .i_c(w_pp_11_09), .ow_sum(w_sum_85), .ow_carry(w_carry_85));
wire w_sum_86, w_carry_86;
math_adder_half HA_86(.i_a(w_pp_12_08), .i_b(w_pp_13_07), .ow_sum(w_sum_86), .ow_carry(w_carry_86));
wire w_sum_87, w_carry_87;
math_adder_carry_save CSA_87(.i_a(w_pp_00_21), .i_b(w_pp_01_20), .i_c(w_pp_02_19), .ow_sum(w_sum_87), .ow_carry(w_carry_87));
wire w_sum_88, w_carry_88;
math_adder_carry_save CSA_88(.i_a(w_pp_03_18), .i_b(w_pp_04_17), .i_c(w_pp_05_16), .ow_sum(w_sum_88), .ow_carry(w_carry_88));
wire w_sum_89, w_carry_89;
math_adder_carry_save CSA_89(.i_a(w_pp_06_15), .i_b(w_pp_07_14), .i_c(w_pp_08_13), .ow_sum(w_sum_89), .ow_carry(w_carry_89));
wire w_sum_90, w_carry_90;
math_adder_carry_save CSA_90(.i_a(w_pp_09_12), .i_b(w_pp_10_11), .i_c(w_pp_11_10), .ow_sum(w_sum_90), .ow_carry(w_carry_90));
wire w_sum_91, w_carry_91;
math_adder_carry_save CSA_91(.i_a(w_pp_12_09), .i_b(w_pp_13_08), .i_c(w_pp_14_07), .ow_sum(w_sum_91), .ow_carry(w_carry_91));
wire w_sum_92, w_carry_92;
math_adder_half HA_92(.i_a(w_pp_15_06), .i_b(w_pp_16_05), .ow_sum(w_sum_92), .ow_carry(w_carry_92));
wire w_sum_93, w_carry_93;
math_adder_carry_save CSA_93(.i_a(w_pp_00_22), .i_b(w_pp_01_21), .i_c(w_pp_02_20), .ow_sum(w_sum_93), .ow_carry(w_carry_93));
wire w_sum_94, w_carry_94;
math_adder_carry_save CSA_94(.i_a(w_pp_03_19), .i_b(w_pp_04_18), .i_c(w_pp_05_17), .ow_sum(w_sum_94), .ow_carry(w_carry_94));
wire w_sum_95, w_carry_95;
math_adder_carry_save CSA_95(.i_a(w_pp_06_16), .i_b(w_pp_07_15), .i_c(w_pp_08_14), .ow_sum(w_sum_95), .ow_carry(w_carry_95));
wire w_sum_96, w_carry_96;
math_adder_carry_save CSA_96(.i_a(w_pp_09_13), .i_b(w_pp_10_12), .i_c(w_pp_11_11), .ow_sum(w_sum_96), .ow_carry(w_carry_96));
wire w_sum_97, w_carry_97;
math_adder_carry_save CSA_97(.i_a(w_pp_12_10), .i_b(w_pp_13_09), .i_c(w_pp_14_08), .ow_sum(w_sum_97), .ow_carry(w_carry_97));
wire w_sum_98, w_carry_98;
math_adder_carry_save CSA_98(.i_a(w_pp_15_07), .i_b(w_pp_16_06), .i_c(w_pp_17_05), .ow_sum(w_sum_98), .ow_carry(w_carry_98));
wire w_sum_99, w_carry_99;
math_adder_half HA_99(.i_a(w_pp_18_04), .i_b(w_pp_19_03), .ow_sum(w_sum_99), .ow_carry(w_carry_99));
wire w_sum_100, w_carry_100;
math_adder_carry_save CSA_100(.i_a(w_pp_00_23), .i_b(w_pp_01_22), .i_c(w_pp_02_21), .ow_sum(w_sum_100), .ow_carry(w_carry_100));
wire w_sum_101, w_carry_101;
math_adder_carry_save CSA_101(.i_a(w_pp_03_20), .i_b(w_pp_04_19), .i_c(w_pp_05_18), .ow_sum(w_sum_101), .ow_carry(w_carry_101));
wire w_sum_102, w_carry_102;
math_adder_carry_save CSA_102(.i_a(w_pp_06_17), .i_b(w_pp_07_16), .i_c(w_pp_08_15), .ow_sum(w_sum_102), .ow_carry(w_carry_102));
wire w_sum_103, w_carry_103;
math_adder_carry_save CSA_103(.i_a(w_pp_09_14), .i_b(w_pp_10_13), .i_c(w_pp_11_12), .ow_sum(w_sum_103), .ow_carry(w_carry_103));
wire w_sum_104, w_carry_104;
math_adder_carry_save CSA_104(.i_a(w_pp_12_11), .i_b(w_pp_13_10), .i_c(w_pp_14_09), .ow_sum(w_sum_104), .ow_carry(w_carry_104));
wire w_sum_105, w_carry_105;
math_adder_carry_save CSA_105(.i_a(w_pp_15_08), .i_b(w_pp_16_07), .i_c(w_pp_17_06), .ow_sum(w_sum_105), .ow_carry(w_carry_105));
wire w_sum_106, w_carry_106;
math_adder_carry_save CSA_106(.i_a(w_pp_18_05), .i_b(w_pp_19_04), .i_c(w_pp_20_03), .ow_sum(w_sum_106), .ow_carry(w_carry_106));
wire w_sum_107, w_carry_107;
math_adder_half HA_107(.i_a(w_pp_21_02), .i_b(w_pp_22_01), .ow_sum(w_sum_107), .ow_carry(w_carry_107));
wire w_sum_108, w_carry_108;
math_adder_carry_save CSA_108(.i_a(w_pp_02_22), .i_b(w_pp_03_21), .i_c(w_pp_04_20), .ow_sum(w_sum_108), .ow_carry(w_carry_108));
wire w_sum_109, w_carry_109;
math_adder_carry_save CSA_109(.i_a(w_pp_05_19), .i_b(w_pp_06_18), .i_c(w_pp_07_17), .ow_sum(w_sum_109), .ow_carry(w_carry_109));
wire w_sum_110, w_carry_110;
math_adder_carry_save CSA_110(.i_a(w_pp_08_16), .i_b(w_pp_09_15), .i_c(w_pp_10_14), .ow_sum(w_sum_110), .ow_carry(w_carry_110));
wire w_sum_111, w_carry_111;
math_adder_carry_save CSA_111(.i_a(w_pp_11_13), .i_b(w_pp_12_12), .i_c(w_pp_13_11), .ow_sum(w_sum_111), .ow_carry(w_carry_111));
wire w_sum_112, w_carry_112;
math_adder_carry_save CSA_112(.i_a(w_pp_14_10), .i_b(w_pp_15_09), .i_c(w_pp_16_08), .ow_sum(w_sum_112), .ow_carry(w_carry_112));
wire w_sum_113, w_carry_113;
math_adder_carry_save CSA_113(.i_a(w_pp_17_07), .i_b(w_pp_18_06), .i_c(w_pp_19_05), .ow_sum(w_sum_113), .ow_carry(w_carry_113));
wire w_sum_114, w_carry_114;
math_adder_carry_save CSA_114(.i_a(w_pp_20_04), .i_b(w_pp_21_03), .i_c(w_pp_22_02), .ow_sum(w_sum_114), .ow_carry(w_carry_114));
wire w_sum_115, w_carry_115;
math_adder_carry_save CSA_115(.i_a(w_pp_23_01), .i_b(w_pp_24_00), .i_c(w_sum_0), .ow_sum(w_sum_115), .ow_carry(w_carry_115));
wire w_sum_116, w_carry_116;
math_adder_carry_save CSA_116(.i_a(w_pp_05_20), .i_b(w_pp_06_19), .i_c(w_pp_07_18), .ow_sum(w_sum_116), .ow_carry(w_carry_116));
wire w_sum_117, w_carry_117;
math_adder_carry_save CSA_117(.i_a(w_pp_08_17), .i_b(w_pp_09_16), .i_c(w_pp_10_15), .ow_sum(w_sum_117), .ow_carry(w_carry_117));
wire w_sum_118, w_carry_118;
math_adder_carry_save CSA_118(.i_a(w_pp_11_14), .i_b(w_pp_12_13), .i_c(w_pp_13_12), .ow_sum(w_sum_118), .ow_carry(w_carry_118));
wire w_sum_119, w_carry_119;
math_adder_carry_save CSA_119(.i_a(w_pp_14_11), .i_b(w_pp_15_10), .i_c(w_pp_16_09), .ow_sum(w_sum_119), .ow_carry(w_carry_119));
wire w_sum_120, w_carry_120;
math_adder_carry_save CSA_120(.i_a(w_pp_17_08), .i_b(w_pp_18_07), .i_c(w_pp_19_06), .ow_sum(w_sum_120), .ow_carry(w_carry_120));
wire w_sum_121, w_carry_121;
math_adder_carry_save CSA_121(.i_a(w_pp_20_05), .i_b(w_pp_21_04), .i_c(w_pp_22_03), .ow_sum(w_sum_121), .ow_carry(w_carry_121));
wire w_sum_122, w_carry_122;
math_adder_carry_save CSA_122(.i_a(w_pp_23_02), .i_b(w_pp_24_01), .i_c(w_pp_25_00), .ow_sum(w_sum_122), .ow_carry(w_carry_122));
wire w_sum_123, w_carry_123;
math_adder_carry_save CSA_123(.i_a(w_carry_0), .i_b(w_sum_1), .i_c(w_sum_2), .ow_sum(w_sum_123), .ow_carry(w_carry_123));
wire w_sum_124, w_carry_124;
math_adder_carry_save CSA_124(.i_a(w_pp_08_18), .i_b(w_pp_09_17), .i_c(w_pp_10_16), .ow_sum(w_sum_124), .ow_carry(w_carry_124));
wire w_sum_125, w_carry_125;
math_adder_carry_save CSA_125(.i_a(w_pp_11_15), .i_b(w_pp_12_14), .i_c(w_pp_13_13), .ow_sum(w_sum_125), .ow_carry(w_carry_125));
wire w_sum_126, w_carry_126;
math_adder_carry_save CSA_126(.i_a(w_pp_14_12), .i_b(w_pp_15_11), .i_c(w_pp_16_10), .ow_sum(w_sum_126), .ow_carry(w_carry_126));
wire w_sum_127, w_carry_127;
math_adder_carry_save CSA_127(.i_a(w_pp_17_09), .i_b(w_pp_18_08), .i_c(w_pp_19_07), .ow_sum(w_sum_127), .ow_carry(w_carry_127));
wire w_sum_128, w_carry_128;
math_adder_carry_save CSA_128(.i_a(w_pp_20_06), .i_b(w_pp_21_05), .i_c(w_pp_22_04), .ow_sum(w_sum_128), .ow_carry(w_carry_128));
wire w_sum_129, w_carry_129;
math_adder_carry_save CSA_129(.i_a(w_pp_23_03), .i_b(w_pp_24_02), .i_c(w_pp_25_01), .ow_sum(w_sum_129), .ow_carry(w_carry_129));
wire w_sum_130, w_carry_130;
math_adder_carry_save CSA_130(.i_a(w_pp_26_00), .i_b(w_carry_1), .i_c(w_carry_2), .ow_sum(w_sum_130), .ow_carry(w_carry_130));
wire w_sum_131, w_carry_131;
math_adder_carry_save CSA_131(.i_a(w_sum_3), .i_b(w_sum_4), .i_c(w_sum_5), .ow_sum(w_sum_131), .ow_carry(w_carry_131));
wire w_sum_132, w_carry_132;
math_adder_carry_save CSA_132(.i_a(w_pp_11_16), .i_b(w_pp_12_15), .i_c(w_pp_13_14), .ow_sum(w_sum_132), .ow_carry(w_carry_132));
wire w_sum_133, w_carry_133;
math_adder_carry_save CSA_133(.i_a(w_pp_14_13), .i_b(w_pp_15_12), .i_c(w_pp_16_11), .ow_sum(w_sum_133), .ow_carry(w_carry_133));
wire w_sum_134, w_carry_134;
math_adder_carry_save CSA_134(.i_a(w_pp_17_10), .i_b(w_pp_18_09), .i_c(w_pp_19_08), .ow_sum(w_sum_134), .ow_carry(w_carry_134));
wire w_sum_135, w_carry_135;
math_adder_carry_save CSA_135(.i_a(w_pp_20_07), .i_b(w_pp_21_06), .i_c(w_pp_22_05), .ow_sum(w_sum_135), .ow_carry(w_carry_135));
wire w_sum_136, w_carry_136;
math_adder_carry_save CSA_136(.i_a(w_pp_23_04), .i_b(w_pp_24_03), .i_c(w_pp_25_02), .ow_sum(w_sum_136), .ow_carry(w_carry_136));
wire w_sum_137, w_carry_137;
math_adder_carry_save CSA_137(.i_a(w_pp_26_01), .i_b(w_pp_27_00), .i_c(w_carry_3), .ow_sum(w_sum_137), .ow_carry(w_carry_137));
wire w_sum_138, w_carry_138;
math_adder_carry_save CSA_138(.i_a(w_carry_4), .i_b(w_carry_5), .i_c(w_sum_6), .ow_sum(w_sum_138), .ow_carry(w_carry_138));
wire w_sum_139, w_carry_139;
math_adder_carry_save CSA_139(.i_a(w_sum_7), .i_b(w_sum_8), .i_c(w_sum_9), .ow_sum(w_sum_139), .ow_carry(w_carry_139));
wire w_sum_140, w_carry_140;
math_adder_carry_save CSA_140(.i_a(w_pp_14_14), .i_b(w_pp_15_13), .i_c(w_pp_16_12), .ow_sum(w_sum_140), .ow_carry(w_carry_140));
wire w_sum_141, w_carry_141;
math_adder_carry_save CSA_141(.i_a(w_pp_17_11), .i_b(w_pp_18_10), .i_c(w_pp_19_09), .ow_sum(w_sum_141), .ow_carry(w_carry_141));
wire w_sum_142, w_carry_142;
math_adder_carry_save CSA_142(.i_a(w_pp_20_08), .i_b(w_pp_21_07), .i_c(w_pp_22_06), .ow_sum(w_sum_142), .ow_carry(w_carry_142));
wire w_sum_143, w_carry_143;
math_adder_carry_save CSA_143(.i_a(w_pp_23_05), .i_b(w_pp_24_04), .i_c(w_pp_25_03), .ow_sum(w_sum_143), .ow_carry(w_carry_143));
wire w_sum_144, w_carry_144;
math_adder_carry_save CSA_144(.i_a(w_pp_26_02), .i_b(w_pp_27_01), .i_c(w_pp_28_00), .ow_sum(w_sum_144), .ow_carry(w_carry_144));
wire w_sum_145, w_carry_145;
math_adder_carry_save CSA_145(.i_a(w_carry_6), .i_b(w_carry_7), .i_c(w_carry_8), .ow_sum(w_sum_145), .ow_carry(w_carry_145));
wire w_sum_146, w_carry_146;
math_adder_carry_save CSA_146(.i_a(w_carry_9), .i_b(w_sum_10), .i_c(w_sum_11), .ow_sum(w_sum_146), .ow_carry(w_carry_146));
wire w_sum_147, w_carry_147;
math_adder_carry_save CSA_147(.i_a(w_sum_12), .i_b(w_sum_13), .i_c(w_sum_14), .ow_sum(w_sum_147), .ow_carry(w_carry_147));
wire w_sum_148, w_carry_148;
math_adder_carry_save CSA_148(.i_a(w_pp_17_12), .i_b(w_pp_18_11), .i_c(w_pp_19_10), .ow_sum(w_sum_148), .ow_carry(w_carry_148));
wire w_sum_149, w_carry_149;
math_adder_carry_save CSA_149(.i_a(w_pp_20_09), .i_b(w_pp_21_08), .i_c(w_pp_22_07), .ow_sum(w_sum_149), .ow_carry(w_carry_149));
wire w_sum_150, w_carry_150;
math_adder_carry_save CSA_150(.i_a(w_pp_23_06), .i_b(w_pp_24_05), .i_c(w_pp_25_04), .ow_sum(w_sum_150), .ow_carry(w_carry_150));
wire w_sum_151, w_carry_151;
math_adder_carry_save CSA_151(.i_a(w_pp_26_03), .i_b(w_pp_27_02), .i_c(w_pp_28_01), .ow_sum(w_sum_151), .ow_carry(w_carry_151));
wire w_sum_152, w_carry_152;
math_adder_carry_save CSA_152(.i_a(w_pp_29_00), .i_b(w_carry_10), .i_c(w_carry_11), .ow_sum(w_sum_152), .ow_carry(w_carry_152));
wire w_sum_153, w_carry_153;
math_adder_carry_save CSA_153(.i_a(w_carry_12), .i_b(w_carry_13), .i_c(w_carry_14), .ow_sum(w_sum_153), .ow_carry(w_carry_153));
wire w_sum_154, w_carry_154;
math_adder_carry_save CSA_154(.i_a(w_sum_15), .i_b(w_sum_16), .i_c(w_sum_17), .ow_sum(w_sum_154), .ow_carry(w_carry_154));
wire w_sum_155, w_carry_155;
math_adder_carry_save CSA_155(.i_a(w_sum_18), .i_b(w_sum_19), .i_c(w_sum_20), .ow_sum(w_sum_155), .ow_carry(w_carry_155));
wire w_sum_156, w_carry_156;
math_adder_carry_save CSA_156(.i_a(w_pp_20_10), .i_b(w_pp_21_09), .i_c(w_pp_22_08), .ow_sum(w_sum_156), .ow_carry(w_carry_156));
wire w_sum_157, w_carry_157;
math_adder_carry_save CSA_157(.i_a(w_pp_23_07), .i_b(w_pp_24_06), .i_c(w_pp_25_05), .ow_sum(w_sum_157), .ow_carry(w_carry_157));
wire w_sum_158, w_carry_158;
math_adder_carry_save CSA_158(.i_a(w_pp_26_04), .i_b(w_pp_27_03), .i_c(w_pp_28_02), .ow_sum(w_sum_158), .ow_carry(w_carry_158));
wire w_sum_159, w_carry_159;
math_adder_carry_save CSA_159(.i_a(w_pp_29_01), .i_b(w_pp_30_00), .i_c(w_carry_15), .ow_sum(w_sum_159), .ow_carry(w_carry_159));
wire w_sum_160, w_carry_160;
math_adder_carry_save CSA_160(.i_a(w_carry_16), .i_b(w_carry_17), .i_c(w_carry_18), .ow_sum(w_sum_160), .ow_carry(w_carry_160));
wire w_sum_161, w_carry_161;
math_adder_carry_save CSA_161(.i_a(w_carry_19), .i_b(w_carry_20), .i_c(w_sum_21), .ow_sum(w_sum_161), .ow_carry(w_carry_161));
wire w_sum_162, w_carry_162;
math_adder_carry_save CSA_162(.i_a(w_sum_22), .i_b(w_sum_23), .i_c(w_sum_24), .ow_sum(w_sum_162), .ow_carry(w_carry_162));
wire w_sum_163, w_carry_163;
math_adder_carry_save CSA_163(.i_a(w_sum_25), .i_b(w_sum_26), .i_c(w_sum_27), .ow_sum(w_sum_163), .ow_carry(w_carry_163));
wire w_sum_164, w_carry_164;
math_adder_carry_save CSA_164(.i_a(w_pp_23_08), .i_b(w_pp_24_07), .i_c(w_pp_25_06), .ow_sum(w_sum_164), .ow_carry(w_carry_164));
wire w_sum_165, w_carry_165;
math_adder_carry_save CSA_165(.i_a(w_pp_26_05), .i_b(w_pp_27_04), .i_c(w_pp_28_03), .ow_sum(w_sum_165), .ow_carry(w_carry_165));
wire w_sum_166, w_carry_166;
math_adder_carry_save CSA_166(.i_a(w_pp_29_02), .i_b(w_pp_30_01), .i_c(w_pp_31_00), .ow_sum(w_sum_166), .ow_carry(w_carry_166));
wire w_sum_167, w_carry_167;
math_adder_carry_save CSA_167(.i_a(w_carry_21), .i_b(w_carry_22), .i_c(w_carry_23), .ow_sum(w_sum_167), .ow_carry(w_carry_167));
wire w_sum_168, w_carry_168;
math_adder_carry_save CSA_168(.i_a(w_carry_24), .i_b(w_carry_25), .i_c(w_carry_26), .ow_sum(w_sum_168), .ow_carry(w_carry_168));
wire w_sum_169, w_carry_169;
math_adder_carry_save CSA_169(.i_a(w_carry_27), .i_b(w_sum_28), .i_c(w_sum_29), .ow_sum(w_sum_169), .ow_carry(w_carry_169));
wire w_sum_170, w_carry_170;
math_adder_carry_save CSA_170(.i_a(w_sum_30), .i_b(w_sum_31), .i_c(w_sum_32), .ow_sum(w_sum_170), .ow_carry(w_carry_170));
wire w_sum_171, w_carry_171;
math_adder_carry_save CSA_171(.i_a(w_sum_33), .i_b(w_sum_34), .i_c(w_sum_35), .ow_sum(w_sum_171), .ow_carry(w_carry_171));
wire w_sum_172, w_carry_172;
math_adder_carry_save CSA_172(.i_a(w_pp_24_08), .i_b(w_pp_25_07), .i_c(w_pp_26_06), .ow_sum(w_sum_172), .ow_carry(w_carry_172));
wire w_sum_173, w_carry_173;
math_adder_carry_save CSA_173(.i_a(w_pp_27_05), .i_b(w_pp_28_04), .i_c(w_pp_29_03), .ow_sum(w_sum_173), .ow_carry(w_carry_173));
wire w_sum_174, w_carry_174;
math_adder_carry_save CSA_174(.i_a(w_pp_30_02), .i_b(w_pp_31_01), .i_c(w_carry_28), .ow_sum(w_sum_174), .ow_carry(w_carry_174));
wire w_sum_175, w_carry_175;
math_adder_carry_save CSA_175(.i_a(w_carry_29), .i_b(w_carry_30), .i_c(w_carry_31), .ow_sum(w_sum_175), .ow_carry(w_carry_175));
wire w_sum_176, w_carry_176;
math_adder_carry_save CSA_176(.i_a(w_carry_32), .i_b(w_carry_33), .i_c(w_carry_34), .ow_sum(w_sum_176), .ow_carry(w_carry_176));
wire w_sum_177, w_carry_177;
math_adder_carry_save CSA_177(.i_a(w_carry_35), .i_b(w_sum_36), .i_c(w_sum_37), .ow_sum(w_sum_177), .ow_carry(w_carry_177));
wire w_sum_178, w_carry_178;
math_adder_carry_save CSA_178(.i_a(w_sum_38), .i_b(w_sum_39), .i_c(w_sum_40), .ow_sum(w_sum_178), .ow_carry(w_carry_178));
wire w_sum_179, w_carry_179;
math_adder_carry_save CSA_179(.i_a(w_sum_41), .i_b(w_sum_42), .i_c(w_sum_43), .ow_sum(w_sum_179), .ow_carry(w_carry_179));
wire w_sum_180, w_carry_180;
math_adder_carry_save CSA_180(.i_a(w_pp_23_10), .i_b(w_pp_24_09), .i_c(w_pp_25_08), .ow_sum(w_sum_180), .ow_carry(w_carry_180));
wire w_sum_181, w_carry_181;
math_adder_carry_save CSA_181(.i_a(w_pp_26_07), .i_b(w_pp_27_06), .i_c(w_pp_28_05), .ow_sum(w_sum_181), .ow_carry(w_carry_181));
wire w_sum_182, w_carry_182;
math_adder_carry_save CSA_182(.i_a(w_pp_29_04), .i_b(w_pp_30_03), .i_c(w_pp_31_02), .ow_sum(w_sum_182), .ow_carry(w_carry_182));
wire w_sum_183, w_carry_183;
math_adder_carry_save CSA_183(.i_a(w_carry_36), .i_b(w_carry_37), .i_c(w_carry_38), .ow_sum(w_sum_183), .ow_carry(w_carry_183));
wire w_sum_184, w_carry_184;
math_adder_carry_save CSA_184(.i_a(w_carry_39), .i_b(w_carry_40), .i_c(w_carry_41), .ow_sum(w_sum_184), .ow_carry(w_carry_184));
wire w_sum_185, w_carry_185;
math_adder_carry_save CSA_185(.i_a(w_carry_42), .i_b(w_carry_43), .i_c(w_sum_44), .ow_sum(w_sum_185), .ow_carry(w_carry_185));
wire w_sum_186, w_carry_186;
math_adder_carry_save CSA_186(.i_a(w_sum_45), .i_b(w_sum_46), .i_c(w_sum_47), .ow_sum(w_sum_186), .ow_carry(w_carry_186));
wire w_sum_187, w_carry_187;
math_adder_carry_save CSA_187(.i_a(w_sum_48), .i_b(w_sum_49), .i_c(w_sum_50), .ow_sum(w_sum_187), .ow_carry(w_carry_187));
wire w_sum_188, w_carry_188;
math_adder_carry_save CSA_188(.i_a(w_pp_21_13), .i_b(w_pp_22_12), .i_c(w_pp_23_11), .ow_sum(w_sum_188), .ow_carry(w_carry_188));
wire w_sum_189, w_carry_189;
math_adder_carry_save CSA_189(.i_a(w_pp_24_10), .i_b(w_pp_25_09), .i_c(w_pp_26_08), .ow_sum(w_sum_189), .ow_carry(w_carry_189));
wire w_sum_190, w_carry_190;
math_adder_carry_save CSA_190(.i_a(w_pp_27_07), .i_b(w_pp_28_06), .i_c(w_pp_29_05), .ow_sum(w_sum_190), .ow_carry(w_carry_190));
wire w_sum_191, w_carry_191;
math_adder_carry_save CSA_191(.i_a(w_pp_30_04), .i_b(w_pp_31_03), .i_c(w_carry_44), .ow_sum(w_sum_191), .ow_carry(w_carry_191));
wire w_sum_192, w_carry_192;
math_adder_carry_save CSA_192(.i_a(w_carry_45), .i_b(w_carry_46), .i_c(w_carry_47), .ow_sum(w_sum_192), .ow_carry(w_carry_192));
wire w_sum_193, w_carry_193;
math_adder_carry_save CSA_193(.i_a(w_carry_48), .i_b(w_carry_49), .i_c(w_carry_50), .ow_sum(w_sum_193), .ow_carry(w_carry_193));
wire w_sum_194, w_carry_194;
math_adder_carry_save CSA_194(.i_a(w_sum_51), .i_b(w_sum_52), .i_c(w_sum_53), .ow_sum(w_sum_194), .ow_carry(w_carry_194));
wire w_sum_195, w_carry_195;
math_adder_carry_save CSA_195(.i_a(w_sum_54), .i_b(w_sum_55), .i_c(w_sum_56), .ow_sum(w_sum_195), .ow_carry(w_carry_195));
wire w_sum_196, w_carry_196;
math_adder_carry_save CSA_196(.i_a(w_pp_19_16), .i_b(w_pp_20_15), .i_c(w_pp_21_14), .ow_sum(w_sum_196), .ow_carry(w_carry_196));
wire w_sum_197, w_carry_197;
math_adder_carry_save CSA_197(.i_a(w_pp_22_13), .i_b(w_pp_23_12), .i_c(w_pp_24_11), .ow_sum(w_sum_197), .ow_carry(w_carry_197));
wire w_sum_198, w_carry_198;
math_adder_carry_save CSA_198(.i_a(w_pp_25_10), .i_b(w_pp_26_09), .i_c(w_pp_27_08), .ow_sum(w_sum_198), .ow_carry(w_carry_198));
wire w_sum_199, w_carry_199;
math_adder_carry_save CSA_199(.i_a(w_pp_28_07), .i_b(w_pp_29_06), .i_c(w_pp_30_05), .ow_sum(w_sum_199), .ow_carry(w_carry_199));
wire w_sum_200, w_carry_200;
math_adder_carry_save CSA_200(.i_a(w_pp_31_04), .i_b(w_carry_51), .i_c(w_carry_52), .ow_sum(w_sum_200), .ow_carry(w_carry_200));
wire w_sum_201, w_carry_201;
math_adder_carry_save CSA_201(.i_a(w_carry_53), .i_b(w_carry_54), .i_c(w_carry_55), .ow_sum(w_sum_201), .ow_carry(w_carry_201));
wire w_sum_202, w_carry_202;
math_adder_carry_save CSA_202(.i_a(w_carry_56), .i_b(w_sum_57), .i_c(w_sum_58), .ow_sum(w_sum_202), .ow_carry(w_carry_202));
wire w_sum_203, w_carry_203;
math_adder_carry_save CSA_203(.i_a(w_sum_59), .i_b(w_sum_60), .i_c(w_sum_61), .ow_sum(w_sum_203), .ow_carry(w_carry_203));
wire w_sum_204, w_carry_204;
math_adder_carry_save CSA_204(.i_a(w_pp_17_19), .i_b(w_pp_18_18), .i_c(w_pp_19_17), .ow_sum(w_sum_204), .ow_carry(w_carry_204));
wire w_sum_205, w_carry_205;
math_adder_carry_save CSA_205(.i_a(w_pp_20_16), .i_b(w_pp_21_15), .i_c(w_pp_22_14), .ow_sum(w_sum_205), .ow_carry(w_carry_205));
wire w_sum_206, w_carry_206;
math_adder_carry_save CSA_206(.i_a(w_pp_23_13), .i_b(w_pp_24_12), .i_c(w_pp_25_11), .ow_sum(w_sum_206), .ow_carry(w_carry_206));
wire w_sum_207, w_carry_207;
math_adder_carry_save CSA_207(.i_a(w_pp_26_10), .i_b(w_pp_27_09), .i_c(w_pp_28_08), .ow_sum(w_sum_207), .ow_carry(w_carry_207));
wire w_sum_208, w_carry_208;
math_adder_carry_save CSA_208(.i_a(w_pp_29_07), .i_b(w_pp_30_06), .i_c(w_pp_31_05), .ow_sum(w_sum_208), .ow_carry(w_carry_208));
wire w_sum_209, w_carry_209;
math_adder_carry_save CSA_209(.i_a(w_carry_57), .i_b(w_carry_58), .i_c(w_carry_59), .ow_sum(w_sum_209), .ow_carry(w_carry_209));
wire w_sum_210, w_carry_210;
math_adder_carry_save CSA_210(.i_a(w_carry_60), .i_b(w_carry_61), .i_c(w_sum_62), .ow_sum(w_sum_210), .ow_carry(w_carry_210));
wire w_sum_211, w_carry_211;
math_adder_carry_save CSA_211(.i_a(w_sum_63), .i_b(w_sum_64), .i_c(w_sum_65), .ow_sum(w_sum_211), .ow_carry(w_carry_211));
wire w_sum_212, w_carry_212;
math_adder_carry_save CSA_212(.i_a(w_pp_15_22), .i_b(w_pp_16_21), .i_c(w_pp_17_20), .ow_sum(w_sum_212), .ow_carry(w_carry_212));
wire w_sum_213, w_carry_213;
math_adder_carry_save CSA_213(.i_a(w_pp_18_19), .i_b(w_pp_19_18), .i_c(w_pp_20_17), .ow_sum(w_sum_213), .ow_carry(w_carry_213));
wire w_sum_214, w_carry_214;
math_adder_carry_save CSA_214(.i_a(w_pp_21_16), .i_b(w_pp_22_15), .i_c(w_pp_23_14), .ow_sum(w_sum_214), .ow_carry(w_carry_214));
wire w_sum_215, w_carry_215;
math_adder_carry_save CSA_215(.i_a(w_pp_24_13), .i_b(w_pp_25_12), .i_c(w_pp_26_11), .ow_sum(w_sum_215), .ow_carry(w_carry_215));
wire w_sum_216, w_carry_216;
math_adder_carry_save CSA_216(.i_a(w_pp_27_10), .i_b(w_pp_28_09), .i_c(w_pp_29_08), .ow_sum(w_sum_216), .ow_carry(w_carry_216));
wire w_sum_217, w_carry_217;
math_adder_carry_save CSA_217(.i_a(w_pp_30_07), .i_b(w_pp_31_06), .i_c(w_carry_62), .ow_sum(w_sum_217), .ow_carry(w_carry_217));
wire w_sum_218, w_carry_218;
math_adder_carry_save CSA_218(.i_a(w_carry_63), .i_b(w_carry_64), .i_c(w_carry_65), .ow_sum(w_sum_218), .ow_carry(w_carry_218));
wire w_sum_219, w_carry_219;
math_adder_carry_save CSA_219(.i_a(w_sum_66), .i_b(w_sum_67), .i_c(w_sum_68), .ow_sum(w_sum_219), .ow_carry(w_carry_219));
wire w_sum_220, w_carry_220;
math_adder_carry_save CSA_220(.i_a(w_pp_13_25), .i_b(w_pp_14_24), .i_c(w_pp_15_23), .ow_sum(w_sum_220), .ow_carry(w_carry_220));
wire w_sum_221, w_carry_221;
math_adder_carry_save CSA_221(.i_a(w_pp_16_22), .i_b(w_pp_17_21), .i_c(w_pp_18_20), .ow_sum(w_sum_221), .ow_carry(w_carry_221));
wire w_sum_222, w_carry_222;
math_adder_carry_save CSA_222(.i_a(w_pp_19_19), .i_b(w_pp_20_18), .i_c(w_pp_21_17), .ow_sum(w_sum_222), .ow_carry(w_carry_222));
wire w_sum_223, w_carry_223;
math_adder_carry_save CSA_223(.i_a(w_pp_22_16), .i_b(w_pp_23_15), .i_c(w_pp_24_14), .ow_sum(w_sum_223), .ow_carry(w_carry_223));
wire w_sum_224, w_carry_224;
math_adder_carry_save CSA_224(.i_a(w_pp_25_13), .i_b(w_pp_26_12), .i_c(w_pp_27_11), .ow_sum(w_sum_224), .ow_carry(w_carry_224));
wire w_sum_225, w_carry_225;
math_adder_carry_save CSA_225(.i_a(w_pp_28_10), .i_b(w_pp_29_09), .i_c(w_pp_30_08), .ow_sum(w_sum_225), .ow_carry(w_carry_225));
wire w_sum_226, w_carry_226;
math_adder_carry_save CSA_226(.i_a(w_pp_31_07), .i_b(w_carry_66), .i_c(w_carry_67), .ow_sum(w_sum_226), .ow_carry(w_carry_226));
wire w_sum_227, w_carry_227;
math_adder_carry_save CSA_227(.i_a(w_carry_68), .i_b(w_sum_69), .i_c(w_sum_70), .ow_sum(w_sum_227), .ow_carry(w_carry_227));
wire w_sum_228, w_carry_228;
math_adder_carry_save CSA_228(.i_a(w_pp_11_28), .i_b(w_pp_12_27), .i_c(w_pp_13_26), .ow_sum(w_sum_228), .ow_carry(w_carry_228));
wire w_sum_229, w_carry_229;
math_adder_carry_save CSA_229(.i_a(w_pp_14_25), .i_b(w_pp_15_24), .i_c(w_pp_16_23), .ow_sum(w_sum_229), .ow_carry(w_carry_229));
wire w_sum_230, w_carry_230;
math_adder_carry_save CSA_230(.i_a(w_pp_17_22), .i_b(w_pp_18_21), .i_c(w_pp_19_20), .ow_sum(w_sum_230), .ow_carry(w_carry_230));
wire w_sum_231, w_carry_231;
math_adder_carry_save CSA_231(.i_a(w_pp_20_19), .i_b(w_pp_21_18), .i_c(w_pp_22_17), .ow_sum(w_sum_231), .ow_carry(w_carry_231));
wire w_sum_232, w_carry_232;
math_adder_carry_save CSA_232(.i_a(w_pp_23_16), .i_b(w_pp_24_15), .i_c(w_pp_25_14), .ow_sum(w_sum_232), .ow_carry(w_carry_232));
wire w_sum_233, w_carry_233;
math_adder_carry_save CSA_233(.i_a(w_pp_26_13), .i_b(w_pp_27_12), .i_c(w_pp_28_11), .ow_sum(w_sum_233), .ow_carry(w_carry_233));
wire w_sum_234, w_carry_234;
math_adder_carry_save CSA_234(.i_a(w_pp_29_10), .i_b(w_pp_30_09), .i_c(w_pp_31_08), .ow_sum(w_sum_234), .ow_carry(w_carry_234));
wire w_sum_235, w_carry_235;
math_adder_carry_save CSA_235(.i_a(w_carry_69), .i_b(w_carry_70), .i_c(w_sum_71), .ow_sum(w_sum_235), .ow_carry(w_carry_235));
wire w_sum_236, w_carry_236;
math_adder_carry_save CSA_236(.i_a(w_pp_09_31), .i_b(w_pp_10_30), .i_c(w_pp_11_29), .ow_sum(w_sum_236), .ow_carry(w_carry_236));
wire w_sum_237, w_carry_237;
math_adder_carry_save CSA_237(.i_a(w_pp_12_28), .i_b(w_pp_13_27), .i_c(w_pp_14_26), .ow_sum(w_sum_237), .ow_carry(w_carry_237));
wire w_sum_238, w_carry_238;
math_adder_carry_save CSA_238(.i_a(w_pp_15_25), .i_b(w_pp_16_24), .i_c(w_pp_17_23), .ow_sum(w_sum_238), .ow_carry(w_carry_238));
wire w_sum_239, w_carry_239;
math_adder_carry_save CSA_239(.i_a(w_pp_18_22), .i_b(w_pp_19_21), .i_c(w_pp_20_20), .ow_sum(w_sum_239), .ow_carry(w_carry_239));
wire w_sum_240, w_carry_240;
math_adder_carry_save CSA_240(.i_a(w_pp_21_19), .i_b(w_pp_22_18), .i_c(w_pp_23_17), .ow_sum(w_sum_240), .ow_carry(w_carry_240));
wire w_sum_241, w_carry_241;
math_adder_carry_save CSA_241(.i_a(w_pp_24_16), .i_b(w_pp_25_15), .i_c(w_pp_26_14), .ow_sum(w_sum_241), .ow_carry(w_carry_241));
wire w_sum_242, w_carry_242;
math_adder_carry_save CSA_242(.i_a(w_pp_27_13), .i_b(w_pp_28_12), .i_c(w_pp_29_11), .ow_sum(w_sum_242), .ow_carry(w_carry_242));
wire w_sum_243, w_carry_243;
math_adder_carry_save CSA_243(.i_a(w_pp_30_10), .i_b(w_pp_31_09), .i_c(w_carry_71), .ow_sum(w_sum_243), .ow_carry(w_carry_243));
wire w_sum_244, w_carry_244;
math_adder_carry_save CSA_244(.i_a(w_pp_10_31), .i_b(w_pp_11_30), .i_c(w_pp_12_29), .ow_sum(w_sum_244), .ow_carry(w_carry_244));
wire w_sum_245, w_carry_245;
math_adder_carry_save CSA_245(.i_a(w_pp_13_28), .i_b(w_pp_14_27), .i_c(w_pp_15_26), .ow_sum(w_sum_245), .ow_carry(w_carry_245));
wire w_sum_246, w_carry_246;
math_adder_carry_save CSA_246(.i_a(w_pp_16_25), .i_b(w_pp_17_24), .i_c(w_pp_18_23), .ow_sum(w_sum_246), .ow_carry(w_carry_246));
wire w_sum_247, w_carry_247;
math_adder_carry_save CSA_247(.i_a(w_pp_19_22), .i_b(w_pp_20_21), .i_c(w_pp_21_20), .ow_sum(w_sum_247), .ow_carry(w_carry_247));
wire w_sum_248, w_carry_248;
math_adder_carry_save CSA_248(.i_a(w_pp_22_19), .i_b(w_pp_23_18), .i_c(w_pp_24_17), .ow_sum(w_sum_248), .ow_carry(w_carry_248));
wire w_sum_249, w_carry_249;
math_adder_carry_save CSA_249(.i_a(w_pp_25_16), .i_b(w_pp_26_15), .i_c(w_pp_27_14), .ow_sum(w_sum_249), .ow_carry(w_carry_249));
wire w_sum_250, w_carry_250;
math_adder_carry_save CSA_250(.i_a(w_pp_28_13), .i_b(w_pp_29_12), .i_c(w_pp_30_11), .ow_sum(w_sum_250), .ow_carry(w_carry_250));
wire w_sum_251, w_carry_251;
math_adder_carry_save CSA_251(.i_a(w_pp_11_31), .i_b(w_pp_12_30), .i_c(w_pp_13_29), .ow_sum(w_sum_251), .ow_carry(w_carry_251));
wire w_sum_252, w_carry_252;
math_adder_carry_save CSA_252(.i_a(w_pp_14_28), .i_b(w_pp_15_27), .i_c(w_pp_16_26), .ow_sum(w_sum_252), .ow_carry(w_carry_252));
wire w_sum_253, w_carry_253;
math_adder_carry_save CSA_253(.i_a(w_pp_17_25), .i_b(w_pp_18_24), .i_c(w_pp_19_23), .ow_sum(w_sum_253), .ow_carry(w_carry_253));
wire w_sum_254, w_carry_254;
math_adder_carry_save CSA_254(.i_a(w_pp_20_22), .i_b(w_pp_21_21), .i_c(w_pp_22_20), .ow_sum(w_sum_254), .ow_carry(w_carry_254));
wire w_sum_255, w_carry_255;
math_adder_carry_save CSA_255(.i_a(w_pp_23_19), .i_b(w_pp_24_18), .i_c(w_pp_25_17), .ow_sum(w_sum_255), .ow_carry(w_carry_255));
wire w_sum_256, w_carry_256;
math_adder_carry_save CSA_256(.i_a(w_pp_26_16), .i_b(w_pp_27_15), .i_c(w_pp_28_14), .ow_sum(w_sum_256), .ow_carry(w_carry_256));
wire w_sum_257, w_carry_257;
math_adder_carry_save CSA_257(.i_a(w_pp_12_31), .i_b(w_pp_13_30), .i_c(w_pp_14_29), .ow_sum(w_sum_257), .ow_carry(w_carry_257));
wire w_sum_258, w_carry_258;
math_adder_carry_save CSA_258(.i_a(w_pp_15_28), .i_b(w_pp_16_27), .i_c(w_pp_17_26), .ow_sum(w_sum_258), .ow_carry(w_carry_258));
wire w_sum_259, w_carry_259;
math_adder_carry_save CSA_259(.i_a(w_pp_18_25), .i_b(w_pp_19_24), .i_c(w_pp_20_23), .ow_sum(w_sum_259), .ow_carry(w_carry_259));
wire w_sum_260, w_carry_260;
math_adder_carry_save CSA_260(.i_a(w_pp_21_22), .i_b(w_pp_22_21), .i_c(w_pp_23_20), .ow_sum(w_sum_260), .ow_carry(w_carry_260));
wire w_sum_261, w_carry_261;
math_adder_carry_save CSA_261(.i_a(w_pp_24_19), .i_b(w_pp_25_18), .i_c(w_pp_26_17), .ow_sum(w_sum_261), .ow_carry(w_carry_261));
wire w_sum_262, w_carry_262;
math_adder_carry_save CSA_262(.i_a(w_pp_13_31), .i_b(w_pp_14_30), .i_c(w_pp_15_29), .ow_sum(w_sum_262), .ow_carry(w_carry_262));
wire w_sum_263, w_carry_263;
math_adder_carry_save CSA_263(.i_a(w_pp_16_28), .i_b(w_pp_17_27), .i_c(w_pp_18_26), .ow_sum(w_sum_263), .ow_carry(w_carry_263));
wire w_sum_264, w_carry_264;
math_adder_carry_save CSA_264(.i_a(w_pp_19_25), .i_b(w_pp_20_24), .i_c(w_pp_21_23), .ow_sum(w_sum_264), .ow_carry(w_carry_264));
wire w_sum_265, w_carry_265;
math_adder_carry_save CSA_265(.i_a(w_pp_22_22), .i_b(w_pp_23_21), .i_c(w_pp_24_20), .ow_sum(w_sum_265), .ow_carry(w_carry_265));
wire w_sum_266, w_carry_266;
math_adder_carry_save CSA_266(.i_a(w_pp_14_31), .i_b(w_pp_15_30), .i_c(w_pp_16_29), .ow_sum(w_sum_266), .ow_carry(w_carry_266));
wire w_sum_267, w_carry_267;
math_adder_carry_save CSA_267(.i_a(w_pp_17_28), .i_b(w_pp_18_27), .i_c(w_pp_19_26), .ow_sum(w_sum_267), .ow_carry(w_carry_267));
wire w_sum_268, w_carry_268;
math_adder_carry_save CSA_268(.i_a(w_pp_20_25), .i_b(w_pp_21_24), .i_c(w_pp_22_23), .ow_sum(w_sum_268), .ow_carry(w_carry_268));
wire w_sum_269, w_carry_269;
math_adder_carry_save CSA_269(.i_a(w_pp_15_31), .i_b(w_pp_16_30), .i_c(w_pp_17_29), .ow_sum(w_sum_269), .ow_carry(w_carry_269));
wire w_sum_270, w_carry_270;
math_adder_carry_save CSA_270(.i_a(w_pp_18_28), .i_b(w_pp_19_27), .i_c(w_pp_20_26), .ow_sum(w_sum_270), .ow_carry(w_carry_270));
wire w_sum_271, w_carry_271;
math_adder_carry_save CSA_271(.i_a(w_pp_16_31), .i_b(w_pp_17_30), .i_c(w_pp_18_29), .ow_sum(w_sum_271), .ow_carry(w_carry_271));
// Stage: 2, Max Height: 12
wire w_sum_272, w_carry_272;
math_adder_half HA_272(.i_a(w_pp_00_12), .i_b(w_pp_01_11), .ow_sum(w_sum_272), .ow_carry(w_carry_272));
wire w_sum_273, w_carry_273;
math_adder_carry_save CSA_273(.i_a(w_pp_00_13), .i_b(w_pp_01_12), .i_c(w_pp_02_11), .ow_sum(w_sum_273), .ow_carry(w_carry_273));
wire w_sum_274, w_carry_274;
math_adder_half HA_274(.i_a(w_pp_03_10), .i_b(w_pp_04_09), .ow_sum(w_sum_274), .ow_carry(w_carry_274));
wire w_sum_275, w_carry_275;
math_adder_carry_save CSA_275(.i_a(w_pp_00_14), .i_b(w_pp_01_13), .i_c(w_pp_02_12), .ow_sum(w_sum_275), .ow_carry(w_carry_275));
wire w_sum_276, w_carry_276;
math_adder_carry_save CSA_276(.i_a(w_pp_03_11), .i_b(w_pp_04_10), .i_c(w_pp_05_09), .ow_sum(w_sum_276), .ow_carry(w_carry_276));
wire w_sum_277, w_carry_277;
math_adder_half HA_277(.i_a(w_pp_06_08), .i_b(w_pp_07_07), .ow_sum(w_sum_277), .ow_carry(w_carry_277));
wire w_sum_278, w_carry_278;
math_adder_carry_save CSA_278(.i_a(w_pp_00_15), .i_b(w_pp_01_14), .i_c(w_pp_02_13), .ow_sum(w_sum_278), .ow_carry(w_carry_278));
wire w_sum_279, w_carry_279;
math_adder_carry_save CSA_279(.i_a(w_pp_03_12), .i_b(w_pp_04_11), .i_c(w_pp_05_10), .ow_sum(w_sum_279), .ow_carry(w_carry_279));
wire w_sum_280, w_carry_280;
math_adder_carry_save CSA_280(.i_a(w_pp_06_09), .i_b(w_pp_07_08), .i_c(w_pp_08_07), .ow_sum(w_sum_280), .ow_carry(w_carry_280));
wire w_sum_281, w_carry_281;
math_adder_half HA_281(.i_a(w_pp_09_06), .i_b(w_pp_10_05), .ow_sum(w_sum_281), .ow_carry(w_carry_281));
wire w_sum_282, w_carry_282;
math_adder_carry_save CSA_282(.i_a(w_pp_02_14), .i_b(w_pp_03_13), .i_c(w_pp_04_12), .ow_sum(w_sum_282), .ow_carry(w_carry_282));
wire w_sum_283, w_carry_283;
math_adder_carry_save CSA_283(.i_a(w_pp_05_11), .i_b(w_pp_06_10), .i_c(w_pp_07_09), .ow_sum(w_sum_283), .ow_carry(w_carry_283));
wire w_sum_284, w_carry_284;
math_adder_carry_save CSA_284(.i_a(w_pp_08_08), .i_b(w_pp_09_07), .i_c(w_pp_10_06), .ow_sum(w_sum_284), .ow_carry(w_carry_284));
wire w_sum_285, w_carry_285;
math_adder_carry_save CSA_285(.i_a(w_pp_11_05), .i_b(w_pp_12_04), .i_c(w_pp_13_03), .ow_sum(w_sum_285), .ow_carry(w_carry_285));
wire w_sum_286, w_carry_286;
math_adder_carry_save CSA_286(.i_a(w_pp_05_12), .i_b(w_pp_06_11), .i_c(w_pp_07_10), .ow_sum(w_sum_286), .ow_carry(w_carry_286));
wire w_sum_287, w_carry_287;
math_adder_carry_save CSA_287(.i_a(w_pp_08_09), .i_b(w_pp_09_08), .i_c(w_pp_10_07), .ow_sum(w_sum_287), .ow_carry(w_carry_287));
wire w_sum_288, w_carry_288;
math_adder_carry_save CSA_288(.i_a(w_pp_11_06), .i_b(w_pp_12_05), .i_c(w_pp_13_04), .ow_sum(w_sum_288), .ow_carry(w_carry_288));
wire w_sum_289, w_carry_289;
math_adder_carry_save CSA_289(.i_a(w_pp_14_03), .i_b(w_pp_15_02), .i_c(w_pp_16_01), .ow_sum(w_sum_289), .ow_carry(w_carry_289));
wire w_sum_290, w_carry_290;
math_adder_carry_save CSA_290(.i_a(w_pp_08_10), .i_b(w_pp_09_09), .i_c(w_pp_10_08), .ow_sum(w_sum_290), .ow_carry(w_carry_290));
wire w_sum_291, w_carry_291;
math_adder_carry_save CSA_291(.i_a(w_pp_11_07), .i_b(w_pp_12_06), .i_c(w_pp_13_05), .ow_sum(w_sum_291), .ow_carry(w_carry_291));
wire w_sum_292, w_carry_292;
math_adder_carry_save CSA_292(.i_a(w_pp_14_04), .i_b(w_pp_15_03), .i_c(w_pp_16_02), .ow_sum(w_sum_292), .ow_carry(w_carry_292));
wire w_sum_293, w_carry_293;
math_adder_carry_save CSA_293(.i_a(w_pp_17_01), .i_b(w_pp_18_00), .i_c(w_carry_73), .ow_sum(w_sum_293), .ow_carry(w_carry_293));
wire w_sum_294, w_carry_294;
math_adder_carry_save CSA_294(.i_a(w_pp_11_08), .i_b(w_pp_12_07), .i_c(w_pp_13_06), .ow_sum(w_sum_294), .ow_carry(w_carry_294));
wire w_sum_295, w_carry_295;
math_adder_carry_save CSA_295(.i_a(w_pp_14_05), .i_b(w_pp_15_04), .i_c(w_pp_16_03), .ow_sum(w_sum_295), .ow_carry(w_carry_295));
wire w_sum_296, w_carry_296;
math_adder_carry_save CSA_296(.i_a(w_pp_17_02), .i_b(w_pp_18_01), .i_c(w_pp_19_00), .ow_sum(w_sum_296), .ow_carry(w_carry_296));
wire w_sum_297, w_carry_297;
math_adder_carry_save CSA_297(.i_a(w_carry_75), .i_b(w_carry_76), .i_c(w_carry_77), .ow_sum(w_sum_297), .ow_carry(w_carry_297));
wire w_sum_298, w_carry_298;
math_adder_carry_save CSA_298(.i_a(w_pp_14_06), .i_b(w_pp_15_05), .i_c(w_pp_16_04), .ow_sum(w_sum_298), .ow_carry(w_carry_298));
wire w_sum_299, w_carry_299;
math_adder_carry_save CSA_299(.i_a(w_pp_17_03), .i_b(w_pp_18_02), .i_c(w_pp_19_01), .ow_sum(w_sum_299), .ow_carry(w_carry_299));
wire w_sum_300, w_carry_300;
math_adder_carry_save CSA_300(.i_a(w_pp_20_00), .i_b(w_carry_78), .i_c(w_carry_79), .ow_sum(w_sum_300), .ow_carry(w_carry_300));
wire w_sum_301, w_carry_301;
math_adder_carry_save CSA_301(.i_a(w_carry_80), .i_b(w_carry_81), .i_c(w_sum_82), .ow_sum(w_sum_301), .ow_carry(w_carry_301));
wire w_sum_302, w_carry_302;
math_adder_carry_save CSA_302(.i_a(w_pp_17_04), .i_b(w_pp_18_03), .i_c(w_pp_19_02), .ow_sum(w_sum_302), .ow_carry(w_carry_302));
wire w_sum_303, w_carry_303;
math_adder_carry_save CSA_303(.i_a(w_pp_20_01), .i_b(w_pp_21_00), .i_c(w_carry_82), .ow_sum(w_sum_303), .ow_carry(w_carry_303));
wire w_sum_304, w_carry_304;
math_adder_carry_save CSA_304(.i_a(w_carry_83), .i_b(w_carry_84), .i_c(w_carry_85), .ow_sum(w_sum_304), .ow_carry(w_carry_304));
wire w_sum_305, w_carry_305;
math_adder_carry_save CSA_305(.i_a(w_carry_86), .i_b(w_sum_87), .i_c(w_sum_88), .ow_sum(w_sum_305), .ow_carry(w_carry_305));
wire w_sum_306, w_carry_306;
math_adder_carry_save CSA_306(.i_a(w_pp_20_02), .i_b(w_pp_21_01), .i_c(w_pp_22_00), .ow_sum(w_sum_306), .ow_carry(w_carry_306));
wire w_sum_307, w_carry_307;
math_adder_carry_save CSA_307(.i_a(w_carry_87), .i_b(w_carry_88), .i_c(w_carry_89), .ow_sum(w_sum_307), .ow_carry(w_carry_307));
wire w_sum_308, w_carry_308;
math_adder_carry_save CSA_308(.i_a(w_carry_90), .i_b(w_carry_91), .i_c(w_carry_92), .ow_sum(w_sum_308), .ow_carry(w_carry_308));
wire w_sum_309, w_carry_309;
math_adder_carry_save CSA_309(.i_a(w_sum_93), .i_b(w_sum_94), .i_c(w_sum_95), .ow_sum(w_sum_309), .ow_carry(w_carry_309));
wire w_sum_310, w_carry_310;
math_adder_carry_save CSA_310(.i_a(w_pp_23_00), .i_b(w_carry_93), .i_c(w_carry_94), .ow_sum(w_sum_310), .ow_carry(w_carry_310));
wire w_sum_311, w_carry_311;
math_adder_carry_save CSA_311(.i_a(w_carry_95), .i_b(w_carry_96), .i_c(w_carry_97), .ow_sum(w_sum_311), .ow_carry(w_carry_311));
wire w_sum_312, w_carry_312;
math_adder_carry_save CSA_312(.i_a(w_carry_98), .i_b(w_carry_99), .i_c(w_sum_100), .ow_sum(w_sum_312), .ow_carry(w_carry_312));
wire w_sum_313, w_carry_313;
math_adder_carry_save CSA_313(.i_a(w_sum_101), .i_b(w_sum_102), .i_c(w_sum_103), .ow_sum(w_sum_313), .ow_carry(w_carry_313));
wire w_sum_314, w_carry_314;
math_adder_carry_save CSA_314(.i_a(w_carry_100), .i_b(w_carry_101), .i_c(w_carry_102), .ow_sum(w_sum_314), .ow_carry(w_carry_314));
wire w_sum_315, w_carry_315;
math_adder_carry_save CSA_315(.i_a(w_carry_103), .i_b(w_carry_104), .i_c(w_carry_105), .ow_sum(w_sum_315), .ow_carry(w_carry_315));
wire w_sum_316, w_carry_316;
math_adder_carry_save CSA_316(.i_a(w_carry_106), .i_b(w_carry_107), .i_c(w_sum_108), .ow_sum(w_sum_316), .ow_carry(w_carry_316));
wire w_sum_317, w_carry_317;
math_adder_carry_save CSA_317(.i_a(w_sum_109), .i_b(w_sum_110), .i_c(w_sum_111), .ow_sum(w_sum_317), .ow_carry(w_carry_317));
wire w_sum_318, w_carry_318;
math_adder_carry_save CSA_318(.i_a(w_carry_108), .i_b(w_carry_109), .i_c(w_carry_110), .ow_sum(w_sum_318), .ow_carry(w_carry_318));
wire w_sum_319, w_carry_319;
math_adder_carry_save CSA_319(.i_a(w_carry_111), .i_b(w_carry_112), .i_c(w_carry_113), .ow_sum(w_sum_319), .ow_carry(w_carry_319));
wire w_sum_320, w_carry_320;
math_adder_carry_save CSA_320(.i_a(w_carry_114), .i_b(w_carry_115), .i_c(w_sum_116), .ow_sum(w_sum_320), .ow_carry(w_carry_320));
wire w_sum_321, w_carry_321;
math_adder_carry_save CSA_321(.i_a(w_sum_117), .i_b(w_sum_118), .i_c(w_sum_119), .ow_sum(w_sum_321), .ow_carry(w_carry_321));
wire w_sum_322, w_carry_322;
math_adder_carry_save CSA_322(.i_a(w_carry_116), .i_b(w_carry_117), .i_c(w_carry_118), .ow_sum(w_sum_322), .ow_carry(w_carry_322));
wire w_sum_323, w_carry_323;
math_adder_carry_save CSA_323(.i_a(w_carry_119), .i_b(w_carry_120), .i_c(w_carry_121), .ow_sum(w_sum_323), .ow_carry(w_carry_323));
wire w_sum_324, w_carry_324;
math_adder_carry_save CSA_324(.i_a(w_carry_122), .i_b(w_carry_123), .i_c(w_sum_124), .ow_sum(w_sum_324), .ow_carry(w_carry_324));
wire w_sum_325, w_carry_325;
math_adder_carry_save CSA_325(.i_a(w_sum_125), .i_b(w_sum_126), .i_c(w_sum_127), .ow_sum(w_sum_325), .ow_carry(w_carry_325));
wire w_sum_326, w_carry_326;
math_adder_carry_save CSA_326(.i_a(w_carry_124), .i_b(w_carry_125), .i_c(w_carry_126), .ow_sum(w_sum_326), .ow_carry(w_carry_326));
wire w_sum_327, w_carry_327;
math_adder_carry_save CSA_327(.i_a(w_carry_127), .i_b(w_carry_128), .i_c(w_carry_129), .ow_sum(w_sum_327), .ow_carry(w_carry_327));
wire w_sum_328, w_carry_328;
math_adder_carry_save CSA_328(.i_a(w_carry_130), .i_b(w_carry_131), .i_c(w_sum_132), .ow_sum(w_sum_328), .ow_carry(w_carry_328));
wire w_sum_329, w_carry_329;
math_adder_carry_save CSA_329(.i_a(w_sum_133), .i_b(w_sum_134), .i_c(w_sum_135), .ow_sum(w_sum_329), .ow_carry(w_carry_329));
wire w_sum_330, w_carry_330;
math_adder_carry_save CSA_330(.i_a(w_carry_132), .i_b(w_carry_133), .i_c(w_carry_134), .ow_sum(w_sum_330), .ow_carry(w_carry_330));
wire w_sum_331, w_carry_331;
math_adder_carry_save CSA_331(.i_a(w_carry_135), .i_b(w_carry_136), .i_c(w_carry_137), .ow_sum(w_sum_331), .ow_carry(w_carry_331));
wire w_sum_332, w_carry_332;
math_adder_carry_save CSA_332(.i_a(w_carry_138), .i_b(w_carry_139), .i_c(w_sum_140), .ow_sum(w_sum_332), .ow_carry(w_carry_332));
wire w_sum_333, w_carry_333;
math_adder_carry_save CSA_333(.i_a(w_sum_141), .i_b(w_sum_142), .i_c(w_sum_143), .ow_sum(w_sum_333), .ow_carry(w_carry_333));
wire w_sum_334, w_carry_334;
math_adder_carry_save CSA_334(.i_a(w_carry_140), .i_b(w_carry_141), .i_c(w_carry_142), .ow_sum(w_sum_334), .ow_carry(w_carry_334));
wire w_sum_335, w_carry_335;
math_adder_carry_save CSA_335(.i_a(w_carry_143), .i_b(w_carry_144), .i_c(w_carry_145), .ow_sum(w_sum_335), .ow_carry(w_carry_335));
wire w_sum_336, w_carry_336;
math_adder_carry_save CSA_336(.i_a(w_carry_146), .i_b(w_carry_147), .i_c(w_sum_148), .ow_sum(w_sum_336), .ow_carry(w_carry_336));
wire w_sum_337, w_carry_337;
math_adder_carry_save CSA_337(.i_a(w_sum_149), .i_b(w_sum_150), .i_c(w_sum_151), .ow_sum(w_sum_337), .ow_carry(w_carry_337));
wire w_sum_338, w_carry_338;
math_adder_carry_save CSA_338(.i_a(w_carry_148), .i_b(w_carry_149), .i_c(w_carry_150), .ow_sum(w_sum_338), .ow_carry(w_carry_338));
wire w_sum_339, w_carry_339;
math_adder_carry_save CSA_339(.i_a(w_carry_151), .i_b(w_carry_152), .i_c(w_carry_153), .ow_sum(w_sum_339), .ow_carry(w_carry_339));
wire w_sum_340, w_carry_340;
math_adder_carry_save CSA_340(.i_a(w_carry_154), .i_b(w_carry_155), .i_c(w_sum_156), .ow_sum(w_sum_340), .ow_carry(w_carry_340));
wire w_sum_341, w_carry_341;
math_adder_carry_save CSA_341(.i_a(w_sum_157), .i_b(w_sum_158), .i_c(w_sum_159), .ow_sum(w_sum_341), .ow_carry(w_carry_341));
wire w_sum_342, w_carry_342;
math_adder_carry_save CSA_342(.i_a(w_carry_156), .i_b(w_carry_157), .i_c(w_carry_158), .ow_sum(w_sum_342), .ow_carry(w_carry_342));
wire w_sum_343, w_carry_343;
math_adder_carry_save CSA_343(.i_a(w_carry_159), .i_b(w_carry_160), .i_c(w_carry_161), .ow_sum(w_sum_343), .ow_carry(w_carry_343));
wire w_sum_344, w_carry_344;
math_adder_carry_save CSA_344(.i_a(w_carry_162), .i_b(w_carry_163), .i_c(w_sum_164), .ow_sum(w_sum_344), .ow_carry(w_carry_344));
wire w_sum_345, w_carry_345;
math_adder_carry_save CSA_345(.i_a(w_sum_165), .i_b(w_sum_166), .i_c(w_sum_167), .ow_sum(w_sum_345), .ow_carry(w_carry_345));
wire w_sum_346, w_carry_346;
math_adder_carry_save CSA_346(.i_a(w_carry_164), .i_b(w_carry_165), .i_c(w_carry_166), .ow_sum(w_sum_346), .ow_carry(w_carry_346));
wire w_sum_347, w_carry_347;
math_adder_carry_save CSA_347(.i_a(w_carry_167), .i_b(w_carry_168), .i_c(w_carry_169), .ow_sum(w_sum_347), .ow_carry(w_carry_347));
wire w_sum_348, w_carry_348;
math_adder_carry_save CSA_348(.i_a(w_carry_170), .i_b(w_carry_171), .i_c(w_sum_172), .ow_sum(w_sum_348), .ow_carry(w_carry_348));
wire w_sum_349, w_carry_349;
math_adder_carry_save CSA_349(.i_a(w_sum_173), .i_b(w_sum_174), .i_c(w_sum_175), .ow_sum(w_sum_349), .ow_carry(w_carry_349));
wire w_sum_350, w_carry_350;
math_adder_carry_save CSA_350(.i_a(w_carry_172), .i_b(w_carry_173), .i_c(w_carry_174), .ow_sum(w_sum_350), .ow_carry(w_carry_350));
wire w_sum_351, w_carry_351;
math_adder_carry_save CSA_351(.i_a(w_carry_175), .i_b(w_carry_176), .i_c(w_carry_177), .ow_sum(w_sum_351), .ow_carry(w_carry_351));
wire w_sum_352, w_carry_352;
math_adder_carry_save CSA_352(.i_a(w_carry_178), .i_b(w_carry_179), .i_c(w_sum_180), .ow_sum(w_sum_352), .ow_carry(w_carry_352));
wire w_sum_353, w_carry_353;
math_adder_carry_save CSA_353(.i_a(w_sum_181), .i_b(w_sum_182), .i_c(w_sum_183), .ow_sum(w_sum_353), .ow_carry(w_carry_353));
wire w_sum_354, w_carry_354;
math_adder_carry_save CSA_354(.i_a(w_carry_180), .i_b(w_carry_181), .i_c(w_carry_182), .ow_sum(w_sum_354), .ow_carry(w_carry_354));
wire w_sum_355, w_carry_355;
math_adder_carry_save CSA_355(.i_a(w_carry_183), .i_b(w_carry_184), .i_c(w_carry_185), .ow_sum(w_sum_355), .ow_carry(w_carry_355));
wire w_sum_356, w_carry_356;
math_adder_carry_save CSA_356(.i_a(w_carry_186), .i_b(w_carry_187), .i_c(w_sum_188), .ow_sum(w_sum_356), .ow_carry(w_carry_356));
wire w_sum_357, w_carry_357;
math_adder_carry_save CSA_357(.i_a(w_sum_189), .i_b(w_sum_190), .i_c(w_sum_191), .ow_sum(w_sum_357), .ow_carry(w_carry_357));
wire w_sum_358, w_carry_358;
math_adder_carry_save CSA_358(.i_a(w_carry_188), .i_b(w_carry_189), .i_c(w_carry_190), .ow_sum(w_sum_358), .ow_carry(w_carry_358));
wire w_sum_359, w_carry_359;
math_adder_carry_save CSA_359(.i_a(w_carry_191), .i_b(w_carry_192), .i_c(w_carry_193), .ow_sum(w_sum_359), .ow_carry(w_carry_359));
wire w_sum_360, w_carry_360;
math_adder_carry_save CSA_360(.i_a(w_carry_194), .i_b(w_carry_195), .i_c(w_sum_196), .ow_sum(w_sum_360), .ow_carry(w_carry_360));
wire w_sum_361, w_carry_361;
math_adder_carry_save CSA_361(.i_a(w_sum_197), .i_b(w_sum_198), .i_c(w_sum_199), .ow_sum(w_sum_361), .ow_carry(w_carry_361));
wire w_sum_362, w_carry_362;
math_adder_carry_save CSA_362(.i_a(w_carry_196), .i_b(w_carry_197), .i_c(w_carry_198), .ow_sum(w_sum_362), .ow_carry(w_carry_362));
wire w_sum_363, w_carry_363;
math_adder_carry_save CSA_363(.i_a(w_carry_199), .i_b(w_carry_200), .i_c(w_carry_201), .ow_sum(w_sum_363), .ow_carry(w_carry_363));
wire w_sum_364, w_carry_364;
math_adder_carry_save CSA_364(.i_a(w_carry_202), .i_b(w_carry_203), .i_c(w_sum_204), .ow_sum(w_sum_364), .ow_carry(w_carry_364));
wire w_sum_365, w_carry_365;
math_adder_carry_save CSA_365(.i_a(w_sum_205), .i_b(w_sum_206), .i_c(w_sum_207), .ow_sum(w_sum_365), .ow_carry(w_carry_365));
wire w_sum_366, w_carry_366;
math_adder_carry_save CSA_366(.i_a(w_carry_204), .i_b(w_carry_205), .i_c(w_carry_206), .ow_sum(w_sum_366), .ow_carry(w_carry_366));
wire w_sum_367, w_carry_367;
math_adder_carry_save CSA_367(.i_a(w_carry_207), .i_b(w_carry_208), .i_c(w_carry_209), .ow_sum(w_sum_367), .ow_carry(w_carry_367));
wire w_sum_368, w_carry_368;
math_adder_carry_save CSA_368(.i_a(w_carry_210), .i_b(w_carry_211), .i_c(w_sum_212), .ow_sum(w_sum_368), .ow_carry(w_carry_368));
wire w_sum_369, w_carry_369;
math_adder_carry_save CSA_369(.i_a(w_sum_213), .i_b(w_sum_214), .i_c(w_sum_215), .ow_sum(w_sum_369), .ow_carry(w_carry_369));
wire w_sum_370, w_carry_370;
math_adder_carry_save CSA_370(.i_a(w_carry_212), .i_b(w_carry_213), .i_c(w_carry_214), .ow_sum(w_sum_370), .ow_carry(w_carry_370));
wire w_sum_371, w_carry_371;
math_adder_carry_save CSA_371(.i_a(w_carry_215), .i_b(w_carry_216), .i_c(w_carry_217), .ow_sum(w_sum_371), .ow_carry(w_carry_371));
wire w_sum_372, w_carry_372;
math_adder_carry_save CSA_372(.i_a(w_carry_218), .i_b(w_carry_219), .i_c(w_sum_220), .ow_sum(w_sum_372), .ow_carry(w_carry_372));
wire w_sum_373, w_carry_373;
math_adder_carry_save CSA_373(.i_a(w_sum_221), .i_b(w_sum_222), .i_c(w_sum_223), .ow_sum(w_sum_373), .ow_carry(w_carry_373));
wire w_sum_374, w_carry_374;
math_adder_carry_save CSA_374(.i_a(w_carry_220), .i_b(w_carry_221), .i_c(w_carry_222), .ow_sum(w_sum_374), .ow_carry(w_carry_374));
wire w_sum_375, w_carry_375;
math_adder_carry_save CSA_375(.i_a(w_carry_223), .i_b(w_carry_224), .i_c(w_carry_225), .ow_sum(w_sum_375), .ow_carry(w_carry_375));
wire w_sum_376, w_carry_376;
math_adder_carry_save CSA_376(.i_a(w_carry_226), .i_b(w_carry_227), .i_c(w_sum_228), .ow_sum(w_sum_376), .ow_carry(w_carry_376));
wire w_sum_377, w_carry_377;
math_adder_carry_save CSA_377(.i_a(w_sum_229), .i_b(w_sum_230), .i_c(w_sum_231), .ow_sum(w_sum_377), .ow_carry(w_carry_377));
wire w_sum_378, w_carry_378;
math_adder_carry_save CSA_378(.i_a(w_carry_228), .i_b(w_carry_229), .i_c(w_carry_230), .ow_sum(w_sum_378), .ow_carry(w_carry_378));
wire w_sum_379, w_carry_379;
math_adder_carry_save CSA_379(.i_a(w_carry_231), .i_b(w_carry_232), .i_c(w_carry_233), .ow_sum(w_sum_379), .ow_carry(w_carry_379));
wire w_sum_380, w_carry_380;
math_adder_carry_save CSA_380(.i_a(w_carry_234), .i_b(w_carry_235), .i_c(w_sum_236), .ow_sum(w_sum_380), .ow_carry(w_carry_380));
wire w_sum_381, w_carry_381;
math_adder_carry_save CSA_381(.i_a(w_sum_237), .i_b(w_sum_238), .i_c(w_sum_239), .ow_sum(w_sum_381), .ow_carry(w_carry_381));
wire w_sum_382, w_carry_382;
math_adder_carry_save CSA_382(.i_a(w_pp_31_10), .i_b(w_carry_236), .i_c(w_carry_237), .ow_sum(w_sum_382), .ow_carry(w_carry_382));
wire w_sum_383, w_carry_383;
math_adder_carry_save CSA_383(.i_a(w_carry_238), .i_b(w_carry_239), .i_c(w_carry_240), .ow_sum(w_sum_383), .ow_carry(w_carry_383));
wire w_sum_384, w_carry_384;
math_adder_carry_save CSA_384(.i_a(w_carry_241), .i_b(w_carry_242), .i_c(w_carry_243), .ow_sum(w_sum_384), .ow_carry(w_carry_384));
wire w_sum_385, w_carry_385;
math_adder_carry_save CSA_385(.i_a(w_sum_244), .i_b(w_sum_245), .i_c(w_sum_246), .ow_sum(w_sum_385), .ow_carry(w_carry_385));
wire w_sum_386, w_carry_386;
math_adder_carry_save CSA_386(.i_a(w_pp_29_13), .i_b(w_pp_30_12), .i_c(w_pp_31_11), .ow_sum(w_sum_386), .ow_carry(w_carry_386));
wire w_sum_387, w_carry_387;
math_adder_carry_save CSA_387(.i_a(w_carry_244), .i_b(w_carry_245), .i_c(w_carry_246), .ow_sum(w_sum_387), .ow_carry(w_carry_387));
wire w_sum_388, w_carry_388;
math_adder_carry_save CSA_388(.i_a(w_carry_247), .i_b(w_carry_248), .i_c(w_carry_249), .ow_sum(w_sum_388), .ow_carry(w_carry_388));
wire w_sum_389, w_carry_389;
math_adder_carry_save CSA_389(.i_a(w_carry_250), .i_b(w_sum_251), .i_c(w_sum_252), .ow_sum(w_sum_389), .ow_carry(w_carry_389));
wire w_sum_390, w_carry_390;
math_adder_carry_save CSA_390(.i_a(w_pp_27_16), .i_b(w_pp_28_15), .i_c(w_pp_29_14), .ow_sum(w_sum_390), .ow_carry(w_carry_390));
wire w_sum_391, w_carry_391;
math_adder_carry_save CSA_391(.i_a(w_pp_30_13), .i_b(w_pp_31_12), .i_c(w_carry_251), .ow_sum(w_sum_391), .ow_carry(w_carry_391));
wire w_sum_392, w_carry_392;
math_adder_carry_save CSA_392(.i_a(w_carry_252), .i_b(w_carry_253), .i_c(w_carry_254), .ow_sum(w_sum_392), .ow_carry(w_carry_392));
wire w_sum_393, w_carry_393;
math_adder_carry_save CSA_393(.i_a(w_carry_255), .i_b(w_carry_256), .i_c(w_sum_257), .ow_sum(w_sum_393), .ow_carry(w_carry_393));
wire w_sum_394, w_carry_394;
math_adder_carry_save CSA_394(.i_a(w_pp_25_19), .i_b(w_pp_26_18), .i_c(w_pp_27_17), .ow_sum(w_sum_394), .ow_carry(w_carry_394));
wire w_sum_395, w_carry_395;
math_adder_carry_save CSA_395(.i_a(w_pp_28_16), .i_b(w_pp_29_15), .i_c(w_pp_30_14), .ow_sum(w_sum_395), .ow_carry(w_carry_395));
wire w_sum_396, w_carry_396;
math_adder_carry_save CSA_396(.i_a(w_pp_31_13), .i_b(w_carry_257), .i_c(w_carry_258), .ow_sum(w_sum_396), .ow_carry(w_carry_396));
wire w_sum_397, w_carry_397;
math_adder_carry_save CSA_397(.i_a(w_carry_259), .i_b(w_carry_260), .i_c(w_carry_261), .ow_sum(w_sum_397), .ow_carry(w_carry_397));
wire w_sum_398, w_carry_398;
math_adder_carry_save CSA_398(.i_a(w_pp_23_22), .i_b(w_pp_24_21), .i_c(w_pp_25_20), .ow_sum(w_sum_398), .ow_carry(w_carry_398));
wire w_sum_399, w_carry_399;
math_adder_carry_save CSA_399(.i_a(w_pp_26_19), .i_b(w_pp_27_18), .i_c(w_pp_28_17), .ow_sum(w_sum_399), .ow_carry(w_carry_399));
wire w_sum_400, w_carry_400;
math_adder_carry_save CSA_400(.i_a(w_pp_29_16), .i_b(w_pp_30_15), .i_c(w_pp_31_14), .ow_sum(w_sum_400), .ow_carry(w_carry_400));
wire w_sum_401, w_carry_401;
math_adder_carry_save CSA_401(.i_a(w_carry_262), .i_b(w_carry_263), .i_c(w_carry_264), .ow_sum(w_sum_401), .ow_carry(w_carry_401));
wire w_sum_402, w_carry_402;
math_adder_carry_save CSA_402(.i_a(w_pp_21_25), .i_b(w_pp_22_24), .i_c(w_pp_23_23), .ow_sum(w_sum_402), .ow_carry(w_carry_402));
wire w_sum_403, w_carry_403;
math_adder_carry_save CSA_403(.i_a(w_pp_24_22), .i_b(w_pp_25_21), .i_c(w_pp_26_20), .ow_sum(w_sum_403), .ow_carry(w_carry_403));
wire w_sum_404, w_carry_404;
math_adder_carry_save CSA_404(.i_a(w_pp_27_19), .i_b(w_pp_28_18), .i_c(w_pp_29_17), .ow_sum(w_sum_404), .ow_carry(w_carry_404));
wire w_sum_405, w_carry_405;
math_adder_carry_save CSA_405(.i_a(w_pp_30_16), .i_b(w_pp_31_15), .i_c(w_carry_266), .ow_sum(w_sum_405), .ow_carry(w_carry_405));
wire w_sum_406, w_carry_406;
math_adder_carry_save CSA_406(.i_a(w_pp_19_28), .i_b(w_pp_20_27), .i_c(w_pp_21_26), .ow_sum(w_sum_406), .ow_carry(w_carry_406));
wire w_sum_407, w_carry_407;
math_adder_carry_save CSA_407(.i_a(w_pp_22_25), .i_b(w_pp_23_24), .i_c(w_pp_24_23), .ow_sum(w_sum_407), .ow_carry(w_carry_407));
wire w_sum_408, w_carry_408;
math_adder_carry_save CSA_408(.i_a(w_pp_25_22), .i_b(w_pp_26_21), .i_c(w_pp_27_20), .ow_sum(w_sum_408), .ow_carry(w_carry_408));
wire w_sum_409, w_carry_409;
math_adder_carry_save CSA_409(.i_a(w_pp_28_19), .i_b(w_pp_29_18), .i_c(w_pp_30_17), .ow_sum(w_sum_409), .ow_carry(w_carry_409));
wire w_sum_410, w_carry_410;
math_adder_carry_save CSA_410(.i_a(w_pp_17_31), .i_b(w_pp_18_30), .i_c(w_pp_19_29), .ow_sum(w_sum_410), .ow_carry(w_carry_410));
wire w_sum_411, w_carry_411;
math_adder_carry_save CSA_411(.i_a(w_pp_20_28), .i_b(w_pp_21_27), .i_c(w_pp_22_26), .ow_sum(w_sum_411), .ow_carry(w_carry_411));
wire w_sum_412, w_carry_412;
math_adder_carry_save CSA_412(.i_a(w_pp_23_25), .i_b(w_pp_24_24), .i_c(w_pp_25_23), .ow_sum(w_sum_412), .ow_carry(w_carry_412));
wire w_sum_413, w_carry_413;
math_adder_carry_save CSA_413(.i_a(w_pp_26_22), .i_b(w_pp_27_21), .i_c(w_pp_28_20), .ow_sum(w_sum_413), .ow_carry(w_carry_413));
wire w_sum_414, w_carry_414;
math_adder_carry_save CSA_414(.i_a(w_pp_18_31), .i_b(w_pp_19_30), .i_c(w_pp_20_29), .ow_sum(w_sum_414), .ow_carry(w_carry_414));
wire w_sum_415, w_carry_415;
math_adder_carry_save CSA_415(.i_a(w_pp_21_28), .i_b(w_pp_22_27), .i_c(w_pp_23_26), .ow_sum(w_sum_415), .ow_carry(w_carry_415));
wire w_sum_416, w_carry_416;
math_adder_carry_save CSA_416(.i_a(w_pp_24_25), .i_b(w_pp_25_24), .i_c(w_pp_26_23), .ow_sum(w_sum_416), .ow_carry(w_carry_416));
wire w_sum_417, w_carry_417;
math_adder_carry_save CSA_417(.i_a(w_pp_19_31), .i_b(w_pp_20_30), .i_c(w_pp_21_29), .ow_sum(w_sum_417), .ow_carry(w_carry_417));
wire w_sum_418, w_carry_418;
math_adder_carry_save CSA_418(.i_a(w_pp_22_28), .i_b(w_pp_23_27), .i_c(w_pp_24_26), .ow_sum(w_sum_418), .ow_carry(w_carry_418));
wire w_sum_419, w_carry_419;
math_adder_carry_save CSA_419(.i_a(w_pp_20_31), .i_b(w_pp_21_30), .i_c(w_pp_22_29), .ow_sum(w_sum_419), .ow_carry(w_carry_419));
// Stage: 3, Max Height: 8
wire w_sum_420, w_carry_420;
math_adder_half HA_420(.i_a(w_pp_00_08), .i_b(w_pp_01_07), .ow_sum(w_sum_420), .ow_carry(w_carry_420));
wire w_sum_421, w_carry_421;
math_adder_carry_save CSA_421(.i_a(w_pp_00_09), .i_b(w_pp_01_08), .i_c(w_pp_02_07), .ow_sum(w_sum_421), .ow_carry(w_carry_421));
wire w_sum_422, w_carry_422;
math_adder_half HA_422(.i_a(w_pp_03_06), .i_b(w_pp_04_05), .ow_sum(w_sum_422), .ow_carry(w_carry_422));
wire w_sum_423, w_carry_423;
math_adder_carry_save CSA_423(.i_a(w_pp_00_10), .i_b(w_pp_01_09), .i_c(w_pp_02_08), .ow_sum(w_sum_423), .ow_carry(w_carry_423));
wire w_sum_424, w_carry_424;
math_adder_carry_save CSA_424(.i_a(w_pp_03_07), .i_b(w_pp_04_06), .i_c(w_pp_05_05), .ow_sum(w_sum_424), .ow_carry(w_carry_424));
wire w_sum_425, w_carry_425;
math_adder_half HA_425(.i_a(w_pp_06_04), .i_b(w_pp_07_03), .ow_sum(w_sum_425), .ow_carry(w_carry_425));
wire w_sum_426, w_carry_426;
math_adder_carry_save CSA_426(.i_a(w_pp_00_11), .i_b(w_pp_01_10), .i_c(w_pp_02_09), .ow_sum(w_sum_426), .ow_carry(w_carry_426));
wire w_sum_427, w_carry_427;
math_adder_carry_save CSA_427(.i_a(w_pp_03_08), .i_b(w_pp_04_07), .i_c(w_pp_05_06), .ow_sum(w_sum_427), .ow_carry(w_carry_427));
wire w_sum_428, w_carry_428;
math_adder_carry_save CSA_428(.i_a(w_pp_06_05), .i_b(w_pp_07_04), .i_c(w_pp_08_03), .ow_sum(w_sum_428), .ow_carry(w_carry_428));
wire w_sum_429, w_carry_429;
math_adder_half HA_429(.i_a(w_pp_09_02), .i_b(w_pp_10_01), .ow_sum(w_sum_429), .ow_carry(w_carry_429));
wire w_sum_430, w_carry_430;
math_adder_carry_save CSA_430(.i_a(w_pp_02_10), .i_b(w_pp_03_09), .i_c(w_pp_04_08), .ow_sum(w_sum_430), .ow_carry(w_carry_430));
wire w_sum_431, w_carry_431;
math_adder_carry_save CSA_431(.i_a(w_pp_05_07), .i_b(w_pp_06_06), .i_c(w_pp_07_05), .ow_sum(w_sum_431), .ow_carry(w_carry_431));
wire w_sum_432, w_carry_432;
math_adder_carry_save CSA_432(.i_a(w_pp_08_04), .i_b(w_pp_09_03), .i_c(w_pp_10_02), .ow_sum(w_sum_432), .ow_carry(w_carry_432));
wire w_sum_433, w_carry_433;
math_adder_carry_save CSA_433(.i_a(w_pp_11_01), .i_b(w_pp_12_00), .i_c(w_sum_272), .ow_sum(w_sum_433), .ow_carry(w_carry_433));
wire w_sum_434, w_carry_434;
math_adder_carry_save CSA_434(.i_a(w_pp_05_08), .i_b(w_pp_06_07), .i_c(w_pp_07_06), .ow_sum(w_sum_434), .ow_carry(w_carry_434));
wire w_sum_435, w_carry_435;
math_adder_carry_save CSA_435(.i_a(w_pp_08_05), .i_b(w_pp_09_04), .i_c(w_pp_10_03), .ow_sum(w_sum_435), .ow_carry(w_carry_435));
wire w_sum_436, w_carry_436;
math_adder_carry_save CSA_436(.i_a(w_pp_11_02), .i_b(w_pp_12_01), .i_c(w_pp_13_00), .ow_sum(w_sum_436), .ow_carry(w_carry_436));
wire w_sum_437, w_carry_437;
math_adder_carry_save CSA_437(.i_a(w_carry_272), .i_b(w_sum_273), .i_c(w_sum_274), .ow_sum(w_sum_437), .ow_carry(w_carry_437));
wire w_sum_438, w_carry_438;
math_adder_carry_save CSA_438(.i_a(w_pp_08_06), .i_b(w_pp_09_05), .i_c(w_pp_10_04), .ow_sum(w_sum_438), .ow_carry(w_carry_438));
wire w_sum_439, w_carry_439;
math_adder_carry_save CSA_439(.i_a(w_pp_11_03), .i_b(w_pp_12_02), .i_c(w_pp_13_01), .ow_sum(w_sum_439), .ow_carry(w_carry_439));
wire w_sum_440, w_carry_440;
math_adder_carry_save CSA_440(.i_a(w_pp_14_00), .i_b(w_carry_273), .i_c(w_carry_274), .ow_sum(w_sum_440), .ow_carry(w_carry_440));
wire w_sum_441, w_carry_441;
math_adder_carry_save CSA_441(.i_a(w_sum_275), .i_b(w_sum_276), .i_c(w_sum_277), .ow_sum(w_sum_441), .ow_carry(w_carry_441));
wire w_sum_442, w_carry_442;
math_adder_carry_save CSA_442(.i_a(w_pp_11_04), .i_b(w_pp_12_03), .i_c(w_pp_13_02), .ow_sum(w_sum_442), .ow_carry(w_carry_442));
wire w_sum_443, w_carry_443;
math_adder_carry_save CSA_443(.i_a(w_pp_14_01), .i_b(w_pp_15_00), .i_c(w_carry_275), .ow_sum(w_sum_443), .ow_carry(w_carry_443));
wire w_sum_444, w_carry_444;
math_adder_carry_save CSA_444(.i_a(w_carry_276), .i_b(w_carry_277), .i_c(w_sum_278), .ow_sum(w_sum_444), .ow_carry(w_carry_444));
wire w_sum_445, w_carry_445;
math_adder_carry_save CSA_445(.i_a(w_sum_279), .i_b(w_sum_280), .i_c(w_sum_281), .ow_sum(w_sum_445), .ow_carry(w_carry_445));
wire w_sum_446, w_carry_446;
math_adder_carry_save CSA_446(.i_a(w_pp_14_02), .i_b(w_pp_15_01), .i_c(w_pp_16_00), .ow_sum(w_sum_446), .ow_carry(w_carry_446));
wire w_sum_447, w_carry_447;
math_adder_carry_save CSA_447(.i_a(w_sum_72), .i_b(w_carry_278), .i_c(w_carry_279), .ow_sum(w_sum_447), .ow_carry(w_carry_447));
wire w_sum_448, w_carry_448;
math_adder_carry_save CSA_448(.i_a(w_carry_280), .i_b(w_carry_281), .i_c(w_sum_282), .ow_sum(w_sum_448), .ow_carry(w_carry_448));
wire w_sum_449, w_carry_449;
math_adder_carry_save CSA_449(.i_a(w_sum_283), .i_b(w_sum_284), .i_c(w_sum_285), .ow_sum(w_sum_449), .ow_carry(w_carry_449));
wire w_sum_450, w_carry_450;
math_adder_carry_save CSA_450(.i_a(w_pp_17_00), .i_b(w_carry_72), .i_c(w_sum_73), .ow_sum(w_sum_450), .ow_carry(w_carry_450));
wire w_sum_451, w_carry_451;
math_adder_carry_save CSA_451(.i_a(w_sum_74), .i_b(w_carry_282), .i_c(w_carry_283), .ow_sum(w_sum_451), .ow_carry(w_carry_451));
wire w_sum_452, w_carry_452;
math_adder_carry_save CSA_452(.i_a(w_carry_284), .i_b(w_carry_285), .i_c(w_sum_286), .ow_sum(w_sum_452), .ow_carry(w_carry_452));
wire w_sum_453, w_carry_453;
math_adder_carry_save CSA_453(.i_a(w_sum_287), .i_b(w_sum_288), .i_c(w_sum_289), .ow_sum(w_sum_453), .ow_carry(w_carry_453));
wire w_sum_454, w_carry_454;
math_adder_carry_save CSA_454(.i_a(w_carry_74), .i_b(w_sum_75), .i_c(w_sum_76), .ow_sum(w_sum_454), .ow_carry(w_carry_454));
wire w_sum_455, w_carry_455;
math_adder_carry_save CSA_455(.i_a(w_sum_77), .i_b(w_carry_286), .i_c(w_carry_287), .ow_sum(w_sum_455), .ow_carry(w_carry_455));
wire w_sum_456, w_carry_456;
math_adder_carry_save CSA_456(.i_a(w_carry_288), .i_b(w_carry_289), .i_c(w_sum_290), .ow_sum(w_sum_456), .ow_carry(w_carry_456));
wire w_sum_457, w_carry_457;
math_adder_carry_save CSA_457(.i_a(w_sum_291), .i_b(w_sum_292), .i_c(w_sum_293), .ow_sum(w_sum_457), .ow_carry(w_carry_457));
wire w_sum_458, w_carry_458;
math_adder_carry_save CSA_458(.i_a(w_sum_78), .i_b(w_sum_79), .i_c(w_sum_80), .ow_sum(w_sum_458), .ow_carry(w_carry_458));
wire w_sum_459, w_carry_459;
math_adder_carry_save CSA_459(.i_a(w_sum_81), .i_b(w_carry_290), .i_c(w_carry_291), .ow_sum(w_sum_459), .ow_carry(w_carry_459));
wire w_sum_460, w_carry_460;
math_adder_carry_save CSA_460(.i_a(w_carry_292), .i_b(w_carry_293), .i_c(w_sum_294), .ow_sum(w_sum_460), .ow_carry(w_carry_460));
wire w_sum_461, w_carry_461;
math_adder_carry_save CSA_461(.i_a(w_sum_295), .i_b(w_sum_296), .i_c(w_sum_297), .ow_sum(w_sum_461), .ow_carry(w_carry_461));
wire w_sum_462, w_carry_462;
math_adder_carry_save CSA_462(.i_a(w_sum_83), .i_b(w_sum_84), .i_c(w_sum_85), .ow_sum(w_sum_462), .ow_carry(w_carry_462));
wire w_sum_463, w_carry_463;
math_adder_carry_save CSA_463(.i_a(w_sum_86), .i_b(w_carry_294), .i_c(w_carry_295), .ow_sum(w_sum_463), .ow_carry(w_carry_463));
wire w_sum_464, w_carry_464;
math_adder_carry_save CSA_464(.i_a(w_carry_296), .i_b(w_carry_297), .i_c(w_sum_298), .ow_sum(w_sum_464), .ow_carry(w_carry_464));
wire w_sum_465, w_carry_465;
math_adder_carry_save CSA_465(.i_a(w_sum_299), .i_b(w_sum_300), .i_c(w_sum_301), .ow_sum(w_sum_465), .ow_carry(w_carry_465));
wire w_sum_466, w_carry_466;
math_adder_carry_save CSA_466(.i_a(w_sum_89), .i_b(w_sum_90), .i_c(w_sum_91), .ow_sum(w_sum_466), .ow_carry(w_carry_466));
wire w_sum_467, w_carry_467;
math_adder_carry_save CSA_467(.i_a(w_sum_92), .i_b(w_carry_298), .i_c(w_carry_299), .ow_sum(w_sum_467), .ow_carry(w_carry_467));
wire w_sum_468, w_carry_468;
math_adder_carry_save CSA_468(.i_a(w_carry_300), .i_b(w_carry_301), .i_c(w_sum_302), .ow_sum(w_sum_468), .ow_carry(w_carry_468));
wire w_sum_469, w_carry_469;
math_adder_carry_save CSA_469(.i_a(w_sum_303), .i_b(w_sum_304), .i_c(w_sum_305), .ow_sum(w_sum_469), .ow_carry(w_carry_469));
wire w_sum_470, w_carry_470;
math_adder_carry_save CSA_470(.i_a(w_sum_96), .i_b(w_sum_97), .i_c(w_sum_98), .ow_sum(w_sum_470), .ow_carry(w_carry_470));
wire w_sum_471, w_carry_471;
math_adder_carry_save CSA_471(.i_a(w_sum_99), .i_b(w_carry_302), .i_c(w_carry_303), .ow_sum(w_sum_471), .ow_carry(w_carry_471));
wire w_sum_472, w_carry_472;
math_adder_carry_save CSA_472(.i_a(w_carry_304), .i_b(w_carry_305), .i_c(w_sum_306), .ow_sum(w_sum_472), .ow_carry(w_carry_472));
wire w_sum_473, w_carry_473;
math_adder_carry_save CSA_473(.i_a(w_sum_307), .i_b(w_sum_308), .i_c(w_sum_309), .ow_sum(w_sum_473), .ow_carry(w_carry_473));
wire w_sum_474, w_carry_474;
math_adder_carry_save CSA_474(.i_a(w_sum_104), .i_b(w_sum_105), .i_c(w_sum_106), .ow_sum(w_sum_474), .ow_carry(w_carry_474));
wire w_sum_475, w_carry_475;
math_adder_carry_save CSA_475(.i_a(w_sum_107), .i_b(w_carry_306), .i_c(w_carry_307), .ow_sum(w_sum_475), .ow_carry(w_carry_475));
wire w_sum_476, w_carry_476;
math_adder_carry_save CSA_476(.i_a(w_carry_308), .i_b(w_carry_309), .i_c(w_sum_310), .ow_sum(w_sum_476), .ow_carry(w_carry_476));
wire w_sum_477, w_carry_477;
math_adder_carry_save CSA_477(.i_a(w_sum_311), .i_b(w_sum_312), .i_c(w_sum_313), .ow_sum(w_sum_477), .ow_carry(w_carry_477));
wire w_sum_478, w_carry_478;
math_adder_carry_save CSA_478(.i_a(w_sum_112), .i_b(w_sum_113), .i_c(w_sum_114), .ow_sum(w_sum_478), .ow_carry(w_carry_478));
wire w_sum_479, w_carry_479;
math_adder_carry_save CSA_479(.i_a(w_sum_115), .i_b(w_carry_310), .i_c(w_carry_311), .ow_sum(w_sum_479), .ow_carry(w_carry_479));
wire w_sum_480, w_carry_480;
math_adder_carry_save CSA_480(.i_a(w_carry_312), .i_b(w_carry_313), .i_c(w_sum_314), .ow_sum(w_sum_480), .ow_carry(w_carry_480));
wire w_sum_481, w_carry_481;
math_adder_carry_save CSA_481(.i_a(w_sum_315), .i_b(w_sum_316), .i_c(w_sum_317), .ow_sum(w_sum_481), .ow_carry(w_carry_481));
wire w_sum_482, w_carry_482;
math_adder_carry_save CSA_482(.i_a(w_sum_120), .i_b(w_sum_121), .i_c(w_sum_122), .ow_sum(w_sum_482), .ow_carry(w_carry_482));
wire w_sum_483, w_carry_483;
math_adder_carry_save CSA_483(.i_a(w_sum_123), .i_b(w_carry_314), .i_c(w_carry_315), .ow_sum(w_sum_483), .ow_carry(w_carry_483));
wire w_sum_484, w_carry_484;
math_adder_carry_save CSA_484(.i_a(w_carry_316), .i_b(w_carry_317), .i_c(w_sum_318), .ow_sum(w_sum_484), .ow_carry(w_carry_484));
wire w_sum_485, w_carry_485;
math_adder_carry_save CSA_485(.i_a(w_sum_319), .i_b(w_sum_320), .i_c(w_sum_321), .ow_sum(w_sum_485), .ow_carry(w_carry_485));
wire w_sum_486, w_carry_486;
math_adder_carry_save CSA_486(.i_a(w_sum_128), .i_b(w_sum_129), .i_c(w_sum_130), .ow_sum(w_sum_486), .ow_carry(w_carry_486));
wire w_sum_487, w_carry_487;
math_adder_carry_save CSA_487(.i_a(w_sum_131), .i_b(w_carry_318), .i_c(w_carry_319), .ow_sum(w_sum_487), .ow_carry(w_carry_487));
wire w_sum_488, w_carry_488;
math_adder_carry_save CSA_488(.i_a(w_carry_320), .i_b(w_carry_321), .i_c(w_sum_322), .ow_sum(w_sum_488), .ow_carry(w_carry_488));
wire w_sum_489, w_carry_489;
math_adder_carry_save CSA_489(.i_a(w_sum_323), .i_b(w_sum_324), .i_c(w_sum_325), .ow_sum(w_sum_489), .ow_carry(w_carry_489));
wire w_sum_490, w_carry_490;
math_adder_carry_save CSA_490(.i_a(w_sum_136), .i_b(w_sum_137), .i_c(w_sum_138), .ow_sum(w_sum_490), .ow_carry(w_carry_490));
wire w_sum_491, w_carry_491;
math_adder_carry_save CSA_491(.i_a(w_sum_139), .i_b(w_carry_322), .i_c(w_carry_323), .ow_sum(w_sum_491), .ow_carry(w_carry_491));
wire w_sum_492, w_carry_492;
math_adder_carry_save CSA_492(.i_a(w_carry_324), .i_b(w_carry_325), .i_c(w_sum_326), .ow_sum(w_sum_492), .ow_carry(w_carry_492));
wire w_sum_493, w_carry_493;
math_adder_carry_save CSA_493(.i_a(w_sum_327), .i_b(w_sum_328), .i_c(w_sum_329), .ow_sum(w_sum_493), .ow_carry(w_carry_493));
wire w_sum_494, w_carry_494;
math_adder_carry_save CSA_494(.i_a(w_sum_144), .i_b(w_sum_145), .i_c(w_sum_146), .ow_sum(w_sum_494), .ow_carry(w_carry_494));
wire w_sum_495, w_carry_495;
math_adder_carry_save CSA_495(.i_a(w_sum_147), .i_b(w_carry_326), .i_c(w_carry_327), .ow_sum(w_sum_495), .ow_carry(w_carry_495));
wire w_sum_496, w_carry_496;
math_adder_carry_save CSA_496(.i_a(w_carry_328), .i_b(w_carry_329), .i_c(w_sum_330), .ow_sum(w_sum_496), .ow_carry(w_carry_496));
wire w_sum_497, w_carry_497;
math_adder_carry_save CSA_497(.i_a(w_sum_331), .i_b(w_sum_332), .i_c(w_sum_333), .ow_sum(w_sum_497), .ow_carry(w_carry_497));
wire w_sum_498, w_carry_498;
math_adder_carry_save CSA_498(.i_a(w_sum_152), .i_b(w_sum_153), .i_c(w_sum_154), .ow_sum(w_sum_498), .ow_carry(w_carry_498));
wire w_sum_499, w_carry_499;
math_adder_carry_save CSA_499(.i_a(w_sum_155), .i_b(w_carry_330), .i_c(w_carry_331), .ow_sum(w_sum_499), .ow_carry(w_carry_499));
wire w_sum_500, w_carry_500;
math_adder_carry_save CSA_500(.i_a(w_carry_332), .i_b(w_carry_333), .i_c(w_sum_334), .ow_sum(w_sum_500), .ow_carry(w_carry_500));
wire w_sum_501, w_carry_501;
math_adder_carry_save CSA_501(.i_a(w_sum_335), .i_b(w_sum_336), .i_c(w_sum_337), .ow_sum(w_sum_501), .ow_carry(w_carry_501));
wire w_sum_502, w_carry_502;
math_adder_carry_save CSA_502(.i_a(w_sum_160), .i_b(w_sum_161), .i_c(w_sum_162), .ow_sum(w_sum_502), .ow_carry(w_carry_502));
wire w_sum_503, w_carry_503;
math_adder_carry_save CSA_503(.i_a(w_sum_163), .i_b(w_carry_334), .i_c(w_carry_335), .ow_sum(w_sum_503), .ow_carry(w_carry_503));
wire w_sum_504, w_carry_504;
math_adder_carry_save CSA_504(.i_a(w_carry_336), .i_b(w_carry_337), .i_c(w_sum_338), .ow_sum(w_sum_504), .ow_carry(w_carry_504));
wire w_sum_505, w_carry_505;
math_adder_carry_save CSA_505(.i_a(w_sum_339), .i_b(w_sum_340), .i_c(w_sum_341), .ow_sum(w_sum_505), .ow_carry(w_carry_505));
wire w_sum_506, w_carry_506;
math_adder_carry_save CSA_506(.i_a(w_sum_168), .i_b(w_sum_169), .i_c(w_sum_170), .ow_sum(w_sum_506), .ow_carry(w_carry_506));
wire w_sum_507, w_carry_507;
math_adder_carry_save CSA_507(.i_a(w_sum_171), .i_b(w_carry_338), .i_c(w_carry_339), .ow_sum(w_sum_507), .ow_carry(w_carry_507));
wire w_sum_508, w_carry_508;
math_adder_carry_save CSA_508(.i_a(w_carry_340), .i_b(w_carry_341), .i_c(w_sum_342), .ow_sum(w_sum_508), .ow_carry(w_carry_508));
wire w_sum_509, w_carry_509;
math_adder_carry_save CSA_509(.i_a(w_sum_343), .i_b(w_sum_344), .i_c(w_sum_345), .ow_sum(w_sum_509), .ow_carry(w_carry_509));
wire w_sum_510, w_carry_510;
math_adder_carry_save CSA_510(.i_a(w_sum_176), .i_b(w_sum_177), .i_c(w_sum_178), .ow_sum(w_sum_510), .ow_carry(w_carry_510));
wire w_sum_511, w_carry_511;
math_adder_carry_save CSA_511(.i_a(w_sum_179), .i_b(w_carry_342), .i_c(w_carry_343), .ow_sum(w_sum_511), .ow_carry(w_carry_511));
wire w_sum_512, w_carry_512;
math_adder_carry_save CSA_512(.i_a(w_carry_344), .i_b(w_carry_345), .i_c(w_sum_346), .ow_sum(w_sum_512), .ow_carry(w_carry_512));
wire w_sum_513, w_carry_513;
math_adder_carry_save CSA_513(.i_a(w_sum_347), .i_b(w_sum_348), .i_c(w_sum_349), .ow_sum(w_sum_513), .ow_carry(w_carry_513));
wire w_sum_514, w_carry_514;
math_adder_carry_save CSA_514(.i_a(w_sum_184), .i_b(w_sum_185), .i_c(w_sum_186), .ow_sum(w_sum_514), .ow_carry(w_carry_514));
wire w_sum_515, w_carry_515;
math_adder_carry_save CSA_515(.i_a(w_sum_187), .i_b(w_carry_346), .i_c(w_carry_347), .ow_sum(w_sum_515), .ow_carry(w_carry_515));
wire w_sum_516, w_carry_516;
math_adder_carry_save CSA_516(.i_a(w_carry_348), .i_b(w_carry_349), .i_c(w_sum_350), .ow_sum(w_sum_516), .ow_carry(w_carry_516));
wire w_sum_517, w_carry_517;
math_adder_carry_save CSA_517(.i_a(w_sum_351), .i_b(w_sum_352), .i_c(w_sum_353), .ow_sum(w_sum_517), .ow_carry(w_carry_517));
wire w_sum_518, w_carry_518;
math_adder_carry_save CSA_518(.i_a(w_sum_192), .i_b(w_sum_193), .i_c(w_sum_194), .ow_sum(w_sum_518), .ow_carry(w_carry_518));
wire w_sum_519, w_carry_519;
math_adder_carry_save CSA_519(.i_a(w_sum_195), .i_b(w_carry_350), .i_c(w_carry_351), .ow_sum(w_sum_519), .ow_carry(w_carry_519));
wire w_sum_520, w_carry_520;
math_adder_carry_save CSA_520(.i_a(w_carry_352), .i_b(w_carry_353), .i_c(w_sum_354), .ow_sum(w_sum_520), .ow_carry(w_carry_520));
wire w_sum_521, w_carry_521;
math_adder_carry_save CSA_521(.i_a(w_sum_355), .i_b(w_sum_356), .i_c(w_sum_357), .ow_sum(w_sum_521), .ow_carry(w_carry_521));
wire w_sum_522, w_carry_522;
math_adder_carry_save CSA_522(.i_a(w_sum_200), .i_b(w_sum_201), .i_c(w_sum_202), .ow_sum(w_sum_522), .ow_carry(w_carry_522));
wire w_sum_523, w_carry_523;
math_adder_carry_save CSA_523(.i_a(w_sum_203), .i_b(w_carry_354), .i_c(w_carry_355), .ow_sum(w_sum_523), .ow_carry(w_carry_523));
wire w_sum_524, w_carry_524;
math_adder_carry_save CSA_524(.i_a(w_carry_356), .i_b(w_carry_357), .i_c(w_sum_358), .ow_sum(w_sum_524), .ow_carry(w_carry_524));
wire w_sum_525, w_carry_525;
math_adder_carry_save CSA_525(.i_a(w_sum_359), .i_b(w_sum_360), .i_c(w_sum_361), .ow_sum(w_sum_525), .ow_carry(w_carry_525));
wire w_sum_526, w_carry_526;
math_adder_carry_save CSA_526(.i_a(w_sum_208), .i_b(w_sum_209), .i_c(w_sum_210), .ow_sum(w_sum_526), .ow_carry(w_carry_526));
wire w_sum_527, w_carry_527;
math_adder_carry_save CSA_527(.i_a(w_sum_211), .i_b(w_carry_358), .i_c(w_carry_359), .ow_sum(w_sum_527), .ow_carry(w_carry_527));
wire w_sum_528, w_carry_528;
math_adder_carry_save CSA_528(.i_a(w_carry_360), .i_b(w_carry_361), .i_c(w_sum_362), .ow_sum(w_sum_528), .ow_carry(w_carry_528));
wire w_sum_529, w_carry_529;
math_adder_carry_save CSA_529(.i_a(w_sum_363), .i_b(w_sum_364), .i_c(w_sum_365), .ow_sum(w_sum_529), .ow_carry(w_carry_529));
wire w_sum_530, w_carry_530;
math_adder_carry_save CSA_530(.i_a(w_sum_216), .i_b(w_sum_217), .i_c(w_sum_218), .ow_sum(w_sum_530), .ow_carry(w_carry_530));
wire w_sum_531, w_carry_531;
math_adder_carry_save CSA_531(.i_a(w_sum_219), .i_b(w_carry_362), .i_c(w_carry_363), .ow_sum(w_sum_531), .ow_carry(w_carry_531));
wire w_sum_532, w_carry_532;
math_adder_carry_save CSA_532(.i_a(w_carry_364), .i_b(w_carry_365), .i_c(w_sum_366), .ow_sum(w_sum_532), .ow_carry(w_carry_532));
wire w_sum_533, w_carry_533;
math_adder_carry_save CSA_533(.i_a(w_sum_367), .i_b(w_sum_368), .i_c(w_sum_369), .ow_sum(w_sum_533), .ow_carry(w_carry_533));
wire w_sum_534, w_carry_534;
math_adder_carry_save CSA_534(.i_a(w_sum_224), .i_b(w_sum_225), .i_c(w_sum_226), .ow_sum(w_sum_534), .ow_carry(w_carry_534));
wire w_sum_535, w_carry_535;
math_adder_carry_save CSA_535(.i_a(w_sum_227), .i_b(w_carry_366), .i_c(w_carry_367), .ow_sum(w_sum_535), .ow_carry(w_carry_535));
wire w_sum_536, w_carry_536;
math_adder_carry_save CSA_536(.i_a(w_carry_368), .i_b(w_carry_369), .i_c(w_sum_370), .ow_sum(w_sum_536), .ow_carry(w_carry_536));
wire w_sum_537, w_carry_537;
math_adder_carry_save CSA_537(.i_a(w_sum_371), .i_b(w_sum_372), .i_c(w_sum_373), .ow_sum(w_sum_537), .ow_carry(w_carry_537));
wire w_sum_538, w_carry_538;
math_adder_carry_save CSA_538(.i_a(w_sum_232), .i_b(w_sum_233), .i_c(w_sum_234), .ow_sum(w_sum_538), .ow_carry(w_carry_538));
wire w_sum_539, w_carry_539;
math_adder_carry_save CSA_539(.i_a(w_sum_235), .i_b(w_carry_370), .i_c(w_carry_371), .ow_sum(w_sum_539), .ow_carry(w_carry_539));
wire w_sum_540, w_carry_540;
math_adder_carry_save CSA_540(.i_a(w_carry_372), .i_b(w_carry_373), .i_c(w_sum_374), .ow_sum(w_sum_540), .ow_carry(w_carry_540));
wire w_sum_541, w_carry_541;
math_adder_carry_save CSA_541(.i_a(w_sum_375), .i_b(w_sum_376), .i_c(w_sum_377), .ow_sum(w_sum_541), .ow_carry(w_carry_541));
wire w_sum_542, w_carry_542;
math_adder_carry_save CSA_542(.i_a(w_sum_240), .i_b(w_sum_241), .i_c(w_sum_242), .ow_sum(w_sum_542), .ow_carry(w_carry_542));
wire w_sum_543, w_carry_543;
math_adder_carry_save CSA_543(.i_a(w_sum_243), .i_b(w_carry_374), .i_c(w_carry_375), .ow_sum(w_sum_543), .ow_carry(w_carry_543));
wire w_sum_544, w_carry_544;
math_adder_carry_save CSA_544(.i_a(w_carry_376), .i_b(w_carry_377), .i_c(w_sum_378), .ow_sum(w_sum_544), .ow_carry(w_carry_544));
wire w_sum_545, w_carry_545;
math_adder_carry_save CSA_545(.i_a(w_sum_379), .i_b(w_sum_380), .i_c(w_sum_381), .ow_sum(w_sum_545), .ow_carry(w_carry_545));
wire w_sum_546, w_carry_546;
math_adder_carry_save CSA_546(.i_a(w_sum_247), .i_b(w_sum_248), .i_c(w_sum_249), .ow_sum(w_sum_546), .ow_carry(w_carry_546));
wire w_sum_547, w_carry_547;
math_adder_carry_save CSA_547(.i_a(w_sum_250), .i_b(w_carry_378), .i_c(w_carry_379), .ow_sum(w_sum_547), .ow_carry(w_carry_547));
wire w_sum_548, w_carry_548;
math_adder_carry_save CSA_548(.i_a(w_carry_380), .i_b(w_carry_381), .i_c(w_sum_382), .ow_sum(w_sum_548), .ow_carry(w_carry_548));
wire w_sum_549, w_carry_549;
math_adder_carry_save CSA_549(.i_a(w_sum_383), .i_b(w_sum_384), .i_c(w_sum_385), .ow_sum(w_sum_549), .ow_carry(w_carry_549));
wire w_sum_550, w_carry_550;
math_adder_carry_save CSA_550(.i_a(w_sum_253), .i_b(w_sum_254), .i_c(w_sum_255), .ow_sum(w_sum_550), .ow_carry(w_carry_550));
wire w_sum_551, w_carry_551;
math_adder_carry_save CSA_551(.i_a(w_sum_256), .i_b(w_carry_382), .i_c(w_carry_383), .ow_sum(w_sum_551), .ow_carry(w_carry_551));
wire w_sum_552, w_carry_552;
math_adder_carry_save CSA_552(.i_a(w_carry_384), .i_b(w_carry_385), .i_c(w_sum_386), .ow_sum(w_sum_552), .ow_carry(w_carry_552));
wire w_sum_553, w_carry_553;
math_adder_carry_save CSA_553(.i_a(w_sum_387), .i_b(w_sum_388), .i_c(w_sum_389), .ow_sum(w_sum_553), .ow_carry(w_carry_553));
wire w_sum_554, w_carry_554;
math_adder_carry_save CSA_554(.i_a(w_sum_258), .i_b(w_sum_259), .i_c(w_sum_260), .ow_sum(w_sum_554), .ow_carry(w_carry_554));
wire w_sum_555, w_carry_555;
math_adder_carry_save CSA_555(.i_a(w_sum_261), .i_b(w_carry_386), .i_c(w_carry_387), .ow_sum(w_sum_555), .ow_carry(w_carry_555));
wire w_sum_556, w_carry_556;
math_adder_carry_save CSA_556(.i_a(w_carry_388), .i_b(w_carry_389), .i_c(w_sum_390), .ow_sum(w_sum_556), .ow_carry(w_carry_556));
wire w_sum_557, w_carry_557;
math_adder_carry_save CSA_557(.i_a(w_sum_391), .i_b(w_sum_392), .i_c(w_sum_393), .ow_sum(w_sum_557), .ow_carry(w_carry_557));
wire w_sum_558, w_carry_558;
math_adder_carry_save CSA_558(.i_a(w_sum_262), .i_b(w_sum_263), .i_c(w_sum_264), .ow_sum(w_sum_558), .ow_carry(w_carry_558));
wire w_sum_559, w_carry_559;
math_adder_carry_save CSA_559(.i_a(w_sum_265), .i_b(w_carry_390), .i_c(w_carry_391), .ow_sum(w_sum_559), .ow_carry(w_carry_559));
wire w_sum_560, w_carry_560;
math_adder_carry_save CSA_560(.i_a(w_carry_392), .i_b(w_carry_393), .i_c(w_sum_394), .ow_sum(w_sum_560), .ow_carry(w_carry_560));
wire w_sum_561, w_carry_561;
math_adder_carry_save CSA_561(.i_a(w_sum_395), .i_b(w_sum_396), .i_c(w_sum_397), .ow_sum(w_sum_561), .ow_carry(w_carry_561));
wire w_sum_562, w_carry_562;
math_adder_carry_save CSA_562(.i_a(w_carry_265), .i_b(w_sum_266), .i_c(w_sum_267), .ow_sum(w_sum_562), .ow_carry(w_carry_562));
wire w_sum_563, w_carry_563;
math_adder_carry_save CSA_563(.i_a(w_sum_268), .i_b(w_carry_394), .i_c(w_carry_395), .ow_sum(w_sum_563), .ow_carry(w_carry_563));
wire w_sum_564, w_carry_564;
math_adder_carry_save CSA_564(.i_a(w_carry_396), .i_b(w_carry_397), .i_c(w_sum_398), .ow_sum(w_sum_564), .ow_carry(w_carry_564));
wire w_sum_565, w_carry_565;
math_adder_carry_save CSA_565(.i_a(w_sum_399), .i_b(w_sum_400), .i_c(w_sum_401), .ow_sum(w_sum_565), .ow_carry(w_carry_565));
wire w_sum_566, w_carry_566;
math_adder_carry_save CSA_566(.i_a(w_carry_267), .i_b(w_carry_268), .i_c(w_sum_269), .ow_sum(w_sum_566), .ow_carry(w_carry_566));
wire w_sum_567, w_carry_567;
math_adder_carry_save CSA_567(.i_a(w_sum_270), .i_b(w_carry_398), .i_c(w_carry_399), .ow_sum(w_sum_567), .ow_carry(w_carry_567));
wire w_sum_568, w_carry_568;
math_adder_carry_save CSA_568(.i_a(w_carry_400), .i_b(w_carry_401), .i_c(w_sum_402), .ow_sum(w_sum_568), .ow_carry(w_carry_568));
wire w_sum_569, w_carry_569;
math_adder_carry_save CSA_569(.i_a(w_sum_403), .i_b(w_sum_404), .i_c(w_sum_405), .ow_sum(w_sum_569), .ow_carry(w_carry_569));
wire w_sum_570, w_carry_570;
math_adder_carry_save CSA_570(.i_a(w_pp_31_16), .i_b(w_carry_269), .i_c(w_carry_270), .ow_sum(w_sum_570), .ow_carry(w_carry_570));
wire w_sum_571, w_carry_571;
math_adder_carry_save CSA_571(.i_a(w_sum_271), .i_b(w_carry_402), .i_c(w_carry_403), .ow_sum(w_sum_571), .ow_carry(w_carry_571));
wire w_sum_572, w_carry_572;
math_adder_carry_save CSA_572(.i_a(w_carry_404), .i_b(w_carry_405), .i_c(w_sum_406), .ow_sum(w_sum_572), .ow_carry(w_carry_572));
wire w_sum_573, w_carry_573;
math_adder_carry_save CSA_573(.i_a(w_sum_407), .i_b(w_sum_408), .i_c(w_sum_409), .ow_sum(w_sum_573), .ow_carry(w_carry_573));
wire w_sum_574, w_carry_574;
math_adder_carry_save CSA_574(.i_a(w_pp_29_19), .i_b(w_pp_30_18), .i_c(w_pp_31_17), .ow_sum(w_sum_574), .ow_carry(w_carry_574));
wire w_sum_575, w_carry_575;
math_adder_carry_save CSA_575(.i_a(w_carry_271), .i_b(w_carry_406), .i_c(w_carry_407), .ow_sum(w_sum_575), .ow_carry(w_carry_575));
wire w_sum_576, w_carry_576;
math_adder_carry_save CSA_576(.i_a(w_carry_408), .i_b(w_carry_409), .i_c(w_sum_410), .ow_sum(w_sum_576), .ow_carry(w_carry_576));
wire w_sum_577, w_carry_577;
math_adder_carry_save CSA_577(.i_a(w_sum_411), .i_b(w_sum_412), .i_c(w_sum_413), .ow_sum(w_sum_577), .ow_carry(w_carry_577));
wire w_sum_578, w_carry_578;
math_adder_carry_save CSA_578(.i_a(w_pp_27_22), .i_b(w_pp_28_21), .i_c(w_pp_29_20), .ow_sum(w_sum_578), .ow_carry(w_carry_578));
wire w_sum_579, w_carry_579;
math_adder_carry_save CSA_579(.i_a(w_pp_30_19), .i_b(w_pp_31_18), .i_c(w_carry_410), .ow_sum(w_sum_579), .ow_carry(w_carry_579));
wire w_sum_580, w_carry_580;
math_adder_carry_save CSA_580(.i_a(w_carry_411), .i_b(w_carry_412), .i_c(w_carry_413), .ow_sum(w_sum_580), .ow_carry(w_carry_580));
wire w_sum_581, w_carry_581;
math_adder_carry_save CSA_581(.i_a(w_sum_414), .i_b(w_sum_415), .i_c(w_sum_416), .ow_sum(w_sum_581), .ow_carry(w_carry_581));
wire w_sum_582, w_carry_582;
math_adder_carry_save CSA_582(.i_a(w_pp_25_25), .i_b(w_pp_26_24), .i_c(w_pp_27_23), .ow_sum(w_sum_582), .ow_carry(w_carry_582));
wire w_sum_583, w_carry_583;
math_adder_carry_save CSA_583(.i_a(w_pp_28_22), .i_b(w_pp_29_21), .i_c(w_pp_30_20), .ow_sum(w_sum_583), .ow_carry(w_carry_583));
wire w_sum_584, w_carry_584;
math_adder_carry_save CSA_584(.i_a(w_pp_31_19), .i_b(w_carry_414), .i_c(w_carry_415), .ow_sum(w_sum_584), .ow_carry(w_carry_584));
wire w_sum_585, w_carry_585;
math_adder_carry_save CSA_585(.i_a(w_carry_416), .i_b(w_sum_417), .i_c(w_sum_418), .ow_sum(w_sum_585), .ow_carry(w_carry_585));
wire w_sum_586, w_carry_586;
math_adder_carry_save CSA_586(.i_a(w_pp_23_28), .i_b(w_pp_24_27), .i_c(w_pp_25_26), .ow_sum(w_sum_586), .ow_carry(w_carry_586));
wire w_sum_587, w_carry_587;
math_adder_carry_save CSA_587(.i_a(w_pp_26_25), .i_b(w_pp_27_24), .i_c(w_pp_28_23), .ow_sum(w_sum_587), .ow_carry(w_carry_587));
wire w_sum_588, w_carry_588;
math_adder_carry_save CSA_588(.i_a(w_pp_29_22), .i_b(w_pp_30_21), .i_c(w_pp_31_20), .ow_sum(w_sum_588), .ow_carry(w_carry_588));
wire w_sum_589, w_carry_589;
math_adder_carry_save CSA_589(.i_a(w_carry_417), .i_b(w_carry_418), .i_c(w_sum_419), .ow_sum(w_sum_589), .ow_carry(w_carry_589));
wire w_sum_590, w_carry_590;
math_adder_carry_save CSA_590(.i_a(w_pp_21_31), .i_b(w_pp_22_30), .i_c(w_pp_23_29), .ow_sum(w_sum_590), .ow_carry(w_carry_590));
wire w_sum_591, w_carry_591;
math_adder_carry_save CSA_591(.i_a(w_pp_24_28), .i_b(w_pp_25_27), .i_c(w_pp_26_26), .ow_sum(w_sum_591), .ow_carry(w_carry_591));
wire w_sum_592, w_carry_592;
math_adder_carry_save CSA_592(.i_a(w_pp_27_25), .i_b(w_pp_28_24), .i_c(w_pp_29_23), .ow_sum(w_sum_592), .ow_carry(w_carry_592));
wire w_sum_593, w_carry_593;
math_adder_carry_save CSA_593(.i_a(w_pp_30_22), .i_b(w_pp_31_21), .i_c(w_carry_419), .ow_sum(w_sum_593), .ow_carry(w_carry_593));
wire w_sum_594, w_carry_594;
math_adder_carry_save CSA_594(.i_a(w_pp_22_31), .i_b(w_pp_23_30), .i_c(w_pp_24_29), .ow_sum(w_sum_594), .ow_carry(w_carry_594));
wire w_sum_595, w_carry_595;
math_adder_carry_save CSA_595(.i_a(w_pp_25_28), .i_b(w_pp_26_27), .i_c(w_pp_27_26), .ow_sum(w_sum_595), .ow_carry(w_carry_595));
wire w_sum_596, w_carry_596;
math_adder_carry_save CSA_596(.i_a(w_pp_28_25), .i_b(w_pp_29_24), .i_c(w_pp_30_23), .ow_sum(w_sum_596), .ow_carry(w_carry_596));
wire w_sum_597, w_carry_597;
math_adder_carry_save CSA_597(.i_a(w_pp_23_31), .i_b(w_pp_24_30), .i_c(w_pp_25_29), .ow_sum(w_sum_597), .ow_carry(w_carry_597));
wire w_sum_598, w_carry_598;
math_adder_carry_save CSA_598(.i_a(w_pp_26_28), .i_b(w_pp_27_27), .i_c(w_pp_28_26), .ow_sum(w_sum_598), .ow_carry(w_carry_598));
wire w_sum_599, w_carry_599;
math_adder_carry_save CSA_599(.i_a(w_pp_24_31), .i_b(w_pp_25_30), .i_c(w_pp_26_29), .ow_sum(w_sum_599), .ow_carry(w_carry_599));
// Stage: 4, Max Height: 6
wire w_sum_600, w_carry_600;
math_adder_half HA_600(.i_a(w_pp_00_06), .i_b(w_pp_01_05), .ow_sum(w_sum_600), .ow_carry(w_carry_600));
wire w_sum_601, w_carry_601;
math_adder_carry_save CSA_601(.i_a(w_pp_00_07), .i_b(w_pp_01_06), .i_c(w_pp_02_05), .ow_sum(w_sum_601), .ow_carry(w_carry_601));
wire w_sum_602, w_carry_602;
math_adder_half HA_602(.i_a(w_pp_03_04), .i_b(w_pp_04_03), .ow_sum(w_sum_602), .ow_carry(w_carry_602));
wire w_sum_603, w_carry_603;
math_adder_carry_save CSA_603(.i_a(w_pp_02_06), .i_b(w_pp_03_05), .i_c(w_pp_04_04), .ow_sum(w_sum_603), .ow_carry(w_carry_603));
wire w_sum_604, w_carry_604;
math_adder_carry_save CSA_604(.i_a(w_pp_05_03), .i_b(w_pp_06_02), .i_c(w_pp_07_01), .ow_sum(w_sum_604), .ow_carry(w_carry_604));
wire w_sum_605, w_carry_605;
math_adder_carry_save CSA_605(.i_a(w_pp_05_04), .i_b(w_pp_06_03), .i_c(w_pp_07_02), .ow_sum(w_sum_605), .ow_carry(w_carry_605));
wire w_sum_606, w_carry_606;
math_adder_carry_save CSA_606(.i_a(w_pp_08_01), .i_b(w_pp_09_00), .i_c(w_carry_420), .ow_sum(w_sum_606), .ow_carry(w_carry_606));
wire w_sum_607, w_carry_607;
math_adder_carry_save CSA_607(.i_a(w_pp_08_02), .i_b(w_pp_09_01), .i_c(w_pp_10_00), .ow_sum(w_sum_607), .ow_carry(w_carry_607));
wire w_sum_608, w_carry_608;
math_adder_carry_save CSA_608(.i_a(w_carry_421), .i_b(w_carry_422), .i_c(w_sum_423), .ow_sum(w_sum_608), .ow_carry(w_carry_608));
wire w_sum_609, w_carry_609;
math_adder_carry_save CSA_609(.i_a(w_pp_11_00), .i_b(w_carry_423), .i_c(w_carry_424), .ow_sum(w_sum_609), .ow_carry(w_carry_609));
wire w_sum_610, w_carry_610;
math_adder_carry_save CSA_610(.i_a(w_carry_425), .i_b(w_sum_426), .i_c(w_sum_427), .ow_sum(w_sum_610), .ow_carry(w_carry_610));
wire w_sum_611, w_carry_611;
math_adder_carry_save CSA_611(.i_a(w_carry_426), .i_b(w_carry_427), .i_c(w_carry_428), .ow_sum(w_sum_611), .ow_carry(w_carry_611));
wire w_sum_612, w_carry_612;
math_adder_carry_save CSA_612(.i_a(w_carry_429), .i_b(w_sum_430), .i_c(w_sum_431), .ow_sum(w_sum_612), .ow_carry(w_carry_612));
wire w_sum_613, w_carry_613;
math_adder_carry_save CSA_613(.i_a(w_carry_430), .i_b(w_carry_431), .i_c(w_carry_432), .ow_sum(w_sum_613), .ow_carry(w_carry_613));
wire w_sum_614, w_carry_614;
math_adder_carry_save CSA_614(.i_a(w_carry_433), .i_b(w_sum_434), .i_c(w_sum_435), .ow_sum(w_sum_614), .ow_carry(w_carry_614));
wire w_sum_615, w_carry_615;
math_adder_carry_save CSA_615(.i_a(w_carry_434), .i_b(w_carry_435), .i_c(w_carry_436), .ow_sum(w_sum_615), .ow_carry(w_carry_615));
wire w_sum_616, w_carry_616;
math_adder_carry_save CSA_616(.i_a(w_carry_437), .i_b(w_sum_438), .i_c(w_sum_439), .ow_sum(w_sum_616), .ow_carry(w_carry_616));
wire w_sum_617, w_carry_617;
math_adder_carry_save CSA_617(.i_a(w_carry_438), .i_b(w_carry_439), .i_c(w_carry_440), .ow_sum(w_sum_617), .ow_carry(w_carry_617));
wire w_sum_618, w_carry_618;
math_adder_carry_save CSA_618(.i_a(w_carry_441), .i_b(w_sum_442), .i_c(w_sum_443), .ow_sum(w_sum_618), .ow_carry(w_carry_618));
wire w_sum_619, w_carry_619;
math_adder_carry_save CSA_619(.i_a(w_carry_442), .i_b(w_carry_443), .i_c(w_carry_444), .ow_sum(w_sum_619), .ow_carry(w_carry_619));
wire w_sum_620, w_carry_620;
math_adder_carry_save CSA_620(.i_a(w_carry_445), .i_b(w_sum_446), .i_c(w_sum_447), .ow_sum(w_sum_620), .ow_carry(w_carry_620));
wire w_sum_621, w_carry_621;
math_adder_carry_save CSA_621(.i_a(w_carry_446), .i_b(w_carry_447), .i_c(w_carry_448), .ow_sum(w_sum_621), .ow_carry(w_carry_621));
wire w_sum_622, w_carry_622;
math_adder_carry_save CSA_622(.i_a(w_carry_449), .i_b(w_sum_450), .i_c(w_sum_451), .ow_sum(w_sum_622), .ow_carry(w_carry_622));
wire w_sum_623, w_carry_623;
math_adder_carry_save CSA_623(.i_a(w_carry_450), .i_b(w_carry_451), .i_c(w_carry_452), .ow_sum(w_sum_623), .ow_carry(w_carry_623));
wire w_sum_624, w_carry_624;
math_adder_carry_save CSA_624(.i_a(w_carry_453), .i_b(w_sum_454), .i_c(w_sum_455), .ow_sum(w_sum_624), .ow_carry(w_carry_624));
wire w_sum_625, w_carry_625;
math_adder_carry_save CSA_625(.i_a(w_carry_454), .i_b(w_carry_455), .i_c(w_carry_456), .ow_sum(w_sum_625), .ow_carry(w_carry_625));
wire w_sum_626, w_carry_626;
math_adder_carry_save CSA_626(.i_a(w_carry_457), .i_b(w_sum_458), .i_c(w_sum_459), .ow_sum(w_sum_626), .ow_carry(w_carry_626));
wire w_sum_627, w_carry_627;
math_adder_carry_save CSA_627(.i_a(w_carry_458), .i_b(w_carry_459), .i_c(w_carry_460), .ow_sum(w_sum_627), .ow_carry(w_carry_627));
wire w_sum_628, w_carry_628;
math_adder_carry_save CSA_628(.i_a(w_carry_461), .i_b(w_sum_462), .i_c(w_sum_463), .ow_sum(w_sum_628), .ow_carry(w_carry_628));
wire w_sum_629, w_carry_629;
math_adder_carry_save CSA_629(.i_a(w_carry_462), .i_b(w_carry_463), .i_c(w_carry_464), .ow_sum(w_sum_629), .ow_carry(w_carry_629));
wire w_sum_630, w_carry_630;
math_adder_carry_save CSA_630(.i_a(w_carry_465), .i_b(w_sum_466), .i_c(w_sum_467), .ow_sum(w_sum_630), .ow_carry(w_carry_630));
wire w_sum_631, w_carry_631;
math_adder_carry_save CSA_631(.i_a(w_carry_466), .i_b(w_carry_467), .i_c(w_carry_468), .ow_sum(w_sum_631), .ow_carry(w_carry_631));
wire w_sum_632, w_carry_632;
math_adder_carry_save CSA_632(.i_a(w_carry_469), .i_b(w_sum_470), .i_c(w_sum_471), .ow_sum(w_sum_632), .ow_carry(w_carry_632));
wire w_sum_633, w_carry_633;
math_adder_carry_save CSA_633(.i_a(w_carry_470), .i_b(w_carry_471), .i_c(w_carry_472), .ow_sum(w_sum_633), .ow_carry(w_carry_633));
wire w_sum_634, w_carry_634;
math_adder_carry_save CSA_634(.i_a(w_carry_473), .i_b(w_sum_474), .i_c(w_sum_475), .ow_sum(w_sum_634), .ow_carry(w_carry_634));
wire w_sum_635, w_carry_635;
math_adder_carry_save CSA_635(.i_a(w_carry_474), .i_b(w_carry_475), .i_c(w_carry_476), .ow_sum(w_sum_635), .ow_carry(w_carry_635));
wire w_sum_636, w_carry_636;
math_adder_carry_save CSA_636(.i_a(w_carry_477), .i_b(w_sum_478), .i_c(w_sum_479), .ow_sum(w_sum_636), .ow_carry(w_carry_636));
wire w_sum_637, w_carry_637;
math_adder_carry_save CSA_637(.i_a(w_carry_478), .i_b(w_carry_479), .i_c(w_carry_480), .ow_sum(w_sum_637), .ow_carry(w_carry_637));
wire w_sum_638, w_carry_638;
math_adder_carry_save CSA_638(.i_a(w_carry_481), .i_b(w_sum_482), .i_c(w_sum_483), .ow_sum(w_sum_638), .ow_carry(w_carry_638));
wire w_sum_639, w_carry_639;
math_adder_carry_save CSA_639(.i_a(w_carry_482), .i_b(w_carry_483), .i_c(w_carry_484), .ow_sum(w_sum_639), .ow_carry(w_carry_639));
wire w_sum_640, w_carry_640;
math_adder_carry_save CSA_640(.i_a(w_carry_485), .i_b(w_sum_486), .i_c(w_sum_487), .ow_sum(w_sum_640), .ow_carry(w_carry_640));
wire w_sum_641, w_carry_641;
math_adder_carry_save CSA_641(.i_a(w_carry_486), .i_b(w_carry_487), .i_c(w_carry_488), .ow_sum(w_sum_641), .ow_carry(w_carry_641));
wire w_sum_642, w_carry_642;
math_adder_carry_save CSA_642(.i_a(w_carry_489), .i_b(w_sum_490), .i_c(w_sum_491), .ow_sum(w_sum_642), .ow_carry(w_carry_642));
wire w_sum_643, w_carry_643;
math_adder_carry_save CSA_643(.i_a(w_carry_490), .i_b(w_carry_491), .i_c(w_carry_492), .ow_sum(w_sum_643), .ow_carry(w_carry_643));
wire w_sum_644, w_carry_644;
math_adder_carry_save CSA_644(.i_a(w_carry_493), .i_b(w_sum_494), .i_c(w_sum_495), .ow_sum(w_sum_644), .ow_carry(w_carry_644));
wire w_sum_645, w_carry_645;
math_adder_carry_save CSA_645(.i_a(w_carry_494), .i_b(w_carry_495), .i_c(w_carry_496), .ow_sum(w_sum_645), .ow_carry(w_carry_645));
wire w_sum_646, w_carry_646;
math_adder_carry_save CSA_646(.i_a(w_carry_497), .i_b(w_sum_498), .i_c(w_sum_499), .ow_sum(w_sum_646), .ow_carry(w_carry_646));
wire w_sum_647, w_carry_647;
math_adder_carry_save CSA_647(.i_a(w_carry_498), .i_b(w_carry_499), .i_c(w_carry_500), .ow_sum(w_sum_647), .ow_carry(w_carry_647));
wire w_sum_648, w_carry_648;
math_adder_carry_save CSA_648(.i_a(w_carry_501), .i_b(w_sum_502), .i_c(w_sum_503), .ow_sum(w_sum_648), .ow_carry(w_carry_648));
wire w_sum_649, w_carry_649;
math_adder_carry_save CSA_649(.i_a(w_carry_502), .i_b(w_carry_503), .i_c(w_carry_504), .ow_sum(w_sum_649), .ow_carry(w_carry_649));
wire w_sum_650, w_carry_650;
math_adder_carry_save CSA_650(.i_a(w_carry_505), .i_b(w_sum_506), .i_c(w_sum_507), .ow_sum(w_sum_650), .ow_carry(w_carry_650));
wire w_sum_651, w_carry_651;
math_adder_carry_save CSA_651(.i_a(w_carry_506), .i_b(w_carry_507), .i_c(w_carry_508), .ow_sum(w_sum_651), .ow_carry(w_carry_651));
wire w_sum_652, w_carry_652;
math_adder_carry_save CSA_652(.i_a(w_carry_509), .i_b(w_sum_510), .i_c(w_sum_511), .ow_sum(w_sum_652), .ow_carry(w_carry_652));
wire w_sum_653, w_carry_653;
math_adder_carry_save CSA_653(.i_a(w_carry_510), .i_b(w_carry_511), .i_c(w_carry_512), .ow_sum(w_sum_653), .ow_carry(w_carry_653));
wire w_sum_654, w_carry_654;
math_adder_carry_save CSA_654(.i_a(w_carry_513), .i_b(w_sum_514), .i_c(w_sum_515), .ow_sum(w_sum_654), .ow_carry(w_carry_654));
wire w_sum_655, w_carry_655;
math_adder_carry_save CSA_655(.i_a(w_carry_514), .i_b(w_carry_515), .i_c(w_carry_516), .ow_sum(w_sum_655), .ow_carry(w_carry_655));
wire w_sum_656, w_carry_656;
math_adder_carry_save CSA_656(.i_a(w_carry_517), .i_b(w_sum_518), .i_c(w_sum_519), .ow_sum(w_sum_656), .ow_carry(w_carry_656));
wire w_sum_657, w_carry_657;
math_adder_carry_save CSA_657(.i_a(w_carry_518), .i_b(w_carry_519), .i_c(w_carry_520), .ow_sum(w_sum_657), .ow_carry(w_carry_657));
wire w_sum_658, w_carry_658;
math_adder_carry_save CSA_658(.i_a(w_carry_521), .i_b(w_sum_522), .i_c(w_sum_523), .ow_sum(w_sum_658), .ow_carry(w_carry_658));
wire w_sum_659, w_carry_659;
math_adder_carry_save CSA_659(.i_a(w_carry_522), .i_b(w_carry_523), .i_c(w_carry_524), .ow_sum(w_sum_659), .ow_carry(w_carry_659));
wire w_sum_660, w_carry_660;
math_adder_carry_save CSA_660(.i_a(w_carry_525), .i_b(w_sum_526), .i_c(w_sum_527), .ow_sum(w_sum_660), .ow_carry(w_carry_660));
wire w_sum_661, w_carry_661;
math_adder_carry_save CSA_661(.i_a(w_carry_526), .i_b(w_carry_527), .i_c(w_carry_528), .ow_sum(w_sum_661), .ow_carry(w_carry_661));
wire w_sum_662, w_carry_662;
math_adder_carry_save CSA_662(.i_a(w_carry_529), .i_b(w_sum_530), .i_c(w_sum_531), .ow_sum(w_sum_662), .ow_carry(w_carry_662));
wire w_sum_663, w_carry_663;
math_adder_carry_save CSA_663(.i_a(w_carry_530), .i_b(w_carry_531), .i_c(w_carry_532), .ow_sum(w_sum_663), .ow_carry(w_carry_663));
wire w_sum_664, w_carry_664;
math_adder_carry_save CSA_664(.i_a(w_carry_533), .i_b(w_sum_534), .i_c(w_sum_535), .ow_sum(w_sum_664), .ow_carry(w_carry_664));
wire w_sum_665, w_carry_665;
math_adder_carry_save CSA_665(.i_a(w_carry_534), .i_b(w_carry_535), .i_c(w_carry_536), .ow_sum(w_sum_665), .ow_carry(w_carry_665));
wire w_sum_666, w_carry_666;
math_adder_carry_save CSA_666(.i_a(w_carry_537), .i_b(w_sum_538), .i_c(w_sum_539), .ow_sum(w_sum_666), .ow_carry(w_carry_666));
wire w_sum_667, w_carry_667;
math_adder_carry_save CSA_667(.i_a(w_carry_538), .i_b(w_carry_539), .i_c(w_carry_540), .ow_sum(w_sum_667), .ow_carry(w_carry_667));
wire w_sum_668, w_carry_668;
math_adder_carry_save CSA_668(.i_a(w_carry_541), .i_b(w_sum_542), .i_c(w_sum_543), .ow_sum(w_sum_668), .ow_carry(w_carry_668));
wire w_sum_669, w_carry_669;
math_adder_carry_save CSA_669(.i_a(w_carry_542), .i_b(w_carry_543), .i_c(w_carry_544), .ow_sum(w_sum_669), .ow_carry(w_carry_669));
wire w_sum_670, w_carry_670;
math_adder_carry_save CSA_670(.i_a(w_carry_545), .i_b(w_sum_546), .i_c(w_sum_547), .ow_sum(w_sum_670), .ow_carry(w_carry_670));
wire w_sum_671, w_carry_671;
math_adder_carry_save CSA_671(.i_a(w_carry_546), .i_b(w_carry_547), .i_c(w_carry_548), .ow_sum(w_sum_671), .ow_carry(w_carry_671));
wire w_sum_672, w_carry_672;
math_adder_carry_save CSA_672(.i_a(w_carry_549), .i_b(w_sum_550), .i_c(w_sum_551), .ow_sum(w_sum_672), .ow_carry(w_carry_672));
wire w_sum_673, w_carry_673;
math_adder_carry_save CSA_673(.i_a(w_carry_550), .i_b(w_carry_551), .i_c(w_carry_552), .ow_sum(w_sum_673), .ow_carry(w_carry_673));
wire w_sum_674, w_carry_674;
math_adder_carry_save CSA_674(.i_a(w_carry_553), .i_b(w_sum_554), .i_c(w_sum_555), .ow_sum(w_sum_674), .ow_carry(w_carry_674));
wire w_sum_675, w_carry_675;
math_adder_carry_save CSA_675(.i_a(w_carry_554), .i_b(w_carry_555), .i_c(w_carry_556), .ow_sum(w_sum_675), .ow_carry(w_carry_675));
wire w_sum_676, w_carry_676;
math_adder_carry_save CSA_676(.i_a(w_carry_557), .i_b(w_sum_558), .i_c(w_sum_559), .ow_sum(w_sum_676), .ow_carry(w_carry_676));
wire w_sum_677, w_carry_677;
math_adder_carry_save CSA_677(.i_a(w_carry_558), .i_b(w_carry_559), .i_c(w_carry_560), .ow_sum(w_sum_677), .ow_carry(w_carry_677));
wire w_sum_678, w_carry_678;
math_adder_carry_save CSA_678(.i_a(w_carry_561), .i_b(w_sum_562), .i_c(w_sum_563), .ow_sum(w_sum_678), .ow_carry(w_carry_678));
wire w_sum_679, w_carry_679;
math_adder_carry_save CSA_679(.i_a(w_carry_562), .i_b(w_carry_563), .i_c(w_carry_564), .ow_sum(w_sum_679), .ow_carry(w_carry_679));
wire w_sum_680, w_carry_680;
math_adder_carry_save CSA_680(.i_a(w_carry_565), .i_b(w_sum_566), .i_c(w_sum_567), .ow_sum(w_sum_680), .ow_carry(w_carry_680));
wire w_sum_681, w_carry_681;
math_adder_carry_save CSA_681(.i_a(w_carry_566), .i_b(w_carry_567), .i_c(w_carry_568), .ow_sum(w_sum_681), .ow_carry(w_carry_681));
wire w_sum_682, w_carry_682;
math_adder_carry_save CSA_682(.i_a(w_carry_569), .i_b(w_sum_570), .i_c(w_sum_571), .ow_sum(w_sum_682), .ow_carry(w_carry_682));
wire w_sum_683, w_carry_683;
math_adder_carry_save CSA_683(.i_a(w_carry_570), .i_b(w_carry_571), .i_c(w_carry_572), .ow_sum(w_sum_683), .ow_carry(w_carry_683));
wire w_sum_684, w_carry_684;
math_adder_carry_save CSA_684(.i_a(w_carry_573), .i_b(w_sum_574), .i_c(w_sum_575), .ow_sum(w_sum_684), .ow_carry(w_carry_684));
wire w_sum_685, w_carry_685;
math_adder_carry_save CSA_685(.i_a(w_carry_574), .i_b(w_carry_575), .i_c(w_carry_576), .ow_sum(w_sum_685), .ow_carry(w_carry_685));
wire w_sum_686, w_carry_686;
math_adder_carry_save CSA_686(.i_a(w_carry_577), .i_b(w_sum_578), .i_c(w_sum_579), .ow_sum(w_sum_686), .ow_carry(w_carry_686));
wire w_sum_687, w_carry_687;
math_adder_carry_save CSA_687(.i_a(w_carry_578), .i_b(w_carry_579), .i_c(w_carry_580), .ow_sum(w_sum_687), .ow_carry(w_carry_687));
wire w_sum_688, w_carry_688;
math_adder_carry_save CSA_688(.i_a(w_carry_581), .i_b(w_sum_582), .i_c(w_sum_583), .ow_sum(w_sum_688), .ow_carry(w_carry_688));
wire w_sum_689, w_carry_689;
math_adder_carry_save CSA_689(.i_a(w_carry_582), .i_b(w_carry_583), .i_c(w_carry_584), .ow_sum(w_sum_689), .ow_carry(w_carry_689));
wire w_sum_690, w_carry_690;
math_adder_carry_save CSA_690(.i_a(w_carry_585), .i_b(w_sum_586), .i_c(w_sum_587), .ow_sum(w_sum_690), .ow_carry(w_carry_690));
wire w_sum_691, w_carry_691;
math_adder_carry_save CSA_691(.i_a(w_carry_586), .i_b(w_carry_587), .i_c(w_carry_588), .ow_sum(w_sum_691), .ow_carry(w_carry_691));
wire w_sum_692, w_carry_692;
math_adder_carry_save CSA_692(.i_a(w_carry_589), .i_b(w_sum_590), .i_c(w_sum_591), .ow_sum(w_sum_692), .ow_carry(w_carry_692));
wire w_sum_693, w_carry_693;
math_adder_carry_save CSA_693(.i_a(w_pp_31_22), .i_b(w_carry_590), .i_c(w_carry_591), .ow_sum(w_sum_693), .ow_carry(w_carry_693));
wire w_sum_694, w_carry_694;
math_adder_carry_save CSA_694(.i_a(w_carry_592), .i_b(w_carry_593), .i_c(w_sum_594), .ow_sum(w_sum_694), .ow_carry(w_carry_694));
wire w_sum_695, w_carry_695;
math_adder_carry_save CSA_695(.i_a(w_pp_29_25), .i_b(w_pp_30_24), .i_c(w_pp_31_23), .ow_sum(w_sum_695), .ow_carry(w_carry_695));
wire w_sum_696, w_carry_696;
math_adder_carry_save CSA_696(.i_a(w_carry_594), .i_b(w_carry_595), .i_c(w_carry_596), .ow_sum(w_sum_696), .ow_carry(w_carry_696));
wire w_sum_697, w_carry_697;
math_adder_carry_save CSA_697(.i_a(w_pp_27_28), .i_b(w_pp_28_27), .i_c(w_pp_29_26), .ow_sum(w_sum_697), .ow_carry(w_carry_697));
wire w_sum_698, w_carry_698;
math_adder_carry_save CSA_698(.i_a(w_pp_30_25), .i_b(w_pp_31_24), .i_c(w_carry_597), .ow_sum(w_sum_698), .ow_carry(w_carry_698));
wire w_sum_699, w_carry_699;
math_adder_carry_save CSA_699(.i_a(w_pp_25_31), .i_b(w_pp_26_30), .i_c(w_pp_27_29), .ow_sum(w_sum_699), .ow_carry(w_carry_699));
wire w_sum_700, w_carry_700;
math_adder_carry_save CSA_700(.i_a(w_pp_28_28), .i_b(w_pp_29_27), .i_c(w_pp_30_26), .ow_sum(w_sum_700), .ow_carry(w_carry_700));
wire w_sum_701, w_carry_701;
math_adder_carry_save CSA_701(.i_a(w_pp_26_31), .i_b(w_pp_27_30), .i_c(w_pp_28_29), .ow_sum(w_sum_701), .ow_carry(w_carry_701));
// Stage: 5, Max Height: 4
wire w_sum_702, w_carry_702;
math_adder_half HA_702(.i_a(w_pp_00_04), .i_b(w_pp_01_03), .ow_sum(w_sum_702), .ow_carry(w_carry_702));
wire w_sum_703, w_carry_703;
math_adder_carry_save CSA_703(.i_a(w_pp_00_05), .i_b(w_pp_01_04), .i_c(w_pp_02_03), .ow_sum(w_sum_703), .ow_carry(w_carry_703));
wire w_sum_704, w_carry_704;
math_adder_half HA_704(.i_a(w_pp_03_02), .i_b(w_pp_04_01), .ow_sum(w_sum_704), .ow_carry(w_carry_704));
wire w_sum_705, w_carry_705;
math_adder_carry_save CSA_705(.i_a(w_pp_02_04), .i_b(w_pp_03_03), .i_c(w_pp_04_02), .ow_sum(w_sum_705), .ow_carry(w_carry_705));
wire w_sum_706, w_carry_706;
math_adder_carry_save CSA_706(.i_a(w_pp_05_01), .i_b(w_pp_06_00), .i_c(w_sum_600), .ow_sum(w_sum_706), .ow_carry(w_carry_706));
wire w_sum_707, w_carry_707;
math_adder_carry_save CSA_707(.i_a(w_pp_05_02), .i_b(w_pp_06_01), .i_c(w_pp_07_00), .ow_sum(w_sum_707), .ow_carry(w_carry_707));
wire w_sum_708, w_carry_708;
math_adder_carry_save CSA_708(.i_a(w_carry_600), .i_b(w_sum_601), .i_c(w_sum_602), .ow_sum(w_sum_708), .ow_carry(w_carry_708));
wire w_sum_709, w_carry_709;
math_adder_carry_save CSA_709(.i_a(w_pp_08_00), .i_b(w_sum_420), .i_c(w_carry_601), .ow_sum(w_sum_709), .ow_carry(w_carry_709));
wire w_sum_710, w_carry_710;
math_adder_carry_save CSA_710(.i_a(w_carry_602), .i_b(w_sum_603), .i_c(w_sum_604), .ow_sum(w_sum_710), .ow_carry(w_carry_710));
wire w_sum_711, w_carry_711;
math_adder_carry_save CSA_711(.i_a(w_sum_421), .i_b(w_sum_422), .i_c(w_carry_603), .ow_sum(w_sum_711), .ow_carry(w_carry_711));
wire w_sum_712, w_carry_712;
math_adder_carry_save CSA_712(.i_a(w_carry_604), .i_b(w_sum_605), .i_c(w_sum_606), .ow_sum(w_sum_712), .ow_carry(w_carry_712));
wire w_sum_713, w_carry_713;
math_adder_carry_save CSA_713(.i_a(w_sum_424), .i_b(w_sum_425), .i_c(w_carry_605), .ow_sum(w_sum_713), .ow_carry(w_carry_713));
wire w_sum_714, w_carry_714;
math_adder_carry_save CSA_714(.i_a(w_carry_606), .i_b(w_sum_607), .i_c(w_sum_608), .ow_sum(w_sum_714), .ow_carry(w_carry_714));
wire w_sum_715, w_carry_715;
math_adder_carry_save CSA_715(.i_a(w_sum_428), .i_b(w_sum_429), .i_c(w_carry_607), .ow_sum(w_sum_715), .ow_carry(w_carry_715));
wire w_sum_716, w_carry_716;
math_adder_carry_save CSA_716(.i_a(w_carry_608), .i_b(w_sum_609), .i_c(w_sum_610), .ow_sum(w_sum_716), .ow_carry(w_carry_716));
wire w_sum_717, w_carry_717;
math_adder_carry_save CSA_717(.i_a(w_sum_432), .i_b(w_sum_433), .i_c(w_carry_609), .ow_sum(w_sum_717), .ow_carry(w_carry_717));
wire w_sum_718, w_carry_718;
math_adder_carry_save CSA_718(.i_a(w_carry_610), .i_b(w_sum_611), .i_c(w_sum_612), .ow_sum(w_sum_718), .ow_carry(w_carry_718));
wire w_sum_719, w_carry_719;
math_adder_carry_save CSA_719(.i_a(w_sum_436), .i_b(w_sum_437), .i_c(w_carry_611), .ow_sum(w_sum_719), .ow_carry(w_carry_719));
wire w_sum_720, w_carry_720;
math_adder_carry_save CSA_720(.i_a(w_carry_612), .i_b(w_sum_613), .i_c(w_sum_614), .ow_sum(w_sum_720), .ow_carry(w_carry_720));
wire w_sum_721, w_carry_721;
math_adder_carry_save CSA_721(.i_a(w_sum_440), .i_b(w_sum_441), .i_c(w_carry_613), .ow_sum(w_sum_721), .ow_carry(w_carry_721));
wire w_sum_722, w_carry_722;
math_adder_carry_save CSA_722(.i_a(w_carry_614), .i_b(w_sum_615), .i_c(w_sum_616), .ow_sum(w_sum_722), .ow_carry(w_carry_722));
wire w_sum_723, w_carry_723;
math_adder_carry_save CSA_723(.i_a(w_sum_444), .i_b(w_sum_445), .i_c(w_carry_615), .ow_sum(w_sum_723), .ow_carry(w_carry_723));
wire w_sum_724, w_carry_724;
math_adder_carry_save CSA_724(.i_a(w_carry_616), .i_b(w_sum_617), .i_c(w_sum_618), .ow_sum(w_sum_724), .ow_carry(w_carry_724));
wire w_sum_725, w_carry_725;
math_adder_carry_save CSA_725(.i_a(w_sum_448), .i_b(w_sum_449), .i_c(w_carry_617), .ow_sum(w_sum_725), .ow_carry(w_carry_725));
wire w_sum_726, w_carry_726;
math_adder_carry_save CSA_726(.i_a(w_carry_618), .i_b(w_sum_619), .i_c(w_sum_620), .ow_sum(w_sum_726), .ow_carry(w_carry_726));
wire w_sum_727, w_carry_727;
math_adder_carry_save CSA_727(.i_a(w_sum_452), .i_b(w_sum_453), .i_c(w_carry_619), .ow_sum(w_sum_727), .ow_carry(w_carry_727));
wire w_sum_728, w_carry_728;
math_adder_carry_save CSA_728(.i_a(w_carry_620), .i_b(w_sum_621), .i_c(w_sum_622), .ow_sum(w_sum_728), .ow_carry(w_carry_728));
wire w_sum_729, w_carry_729;
math_adder_carry_save CSA_729(.i_a(w_sum_456), .i_b(w_sum_457), .i_c(w_carry_621), .ow_sum(w_sum_729), .ow_carry(w_carry_729));
wire w_sum_730, w_carry_730;
math_adder_carry_save CSA_730(.i_a(w_carry_622), .i_b(w_sum_623), .i_c(w_sum_624), .ow_sum(w_sum_730), .ow_carry(w_carry_730));
wire w_sum_731, w_carry_731;
math_adder_carry_save CSA_731(.i_a(w_sum_460), .i_b(w_sum_461), .i_c(w_carry_623), .ow_sum(w_sum_731), .ow_carry(w_carry_731));
wire w_sum_732, w_carry_732;
math_adder_carry_save CSA_732(.i_a(w_carry_624), .i_b(w_sum_625), .i_c(w_sum_626), .ow_sum(w_sum_732), .ow_carry(w_carry_732));
wire w_sum_733, w_carry_733;
math_adder_carry_save CSA_733(.i_a(w_sum_464), .i_b(w_sum_465), .i_c(w_carry_625), .ow_sum(w_sum_733), .ow_carry(w_carry_733));
wire w_sum_734, w_carry_734;
math_adder_carry_save CSA_734(.i_a(w_carry_626), .i_b(w_sum_627), .i_c(w_sum_628), .ow_sum(w_sum_734), .ow_carry(w_carry_734));
wire w_sum_735, w_carry_735;
math_adder_carry_save CSA_735(.i_a(w_sum_468), .i_b(w_sum_469), .i_c(w_carry_627), .ow_sum(w_sum_735), .ow_carry(w_carry_735));
wire w_sum_736, w_carry_736;
math_adder_carry_save CSA_736(.i_a(w_carry_628), .i_b(w_sum_629), .i_c(w_sum_630), .ow_sum(w_sum_736), .ow_carry(w_carry_736));
wire w_sum_737, w_carry_737;
math_adder_carry_save CSA_737(.i_a(w_sum_472), .i_b(w_sum_473), .i_c(w_carry_629), .ow_sum(w_sum_737), .ow_carry(w_carry_737));
wire w_sum_738, w_carry_738;
math_adder_carry_save CSA_738(.i_a(w_carry_630), .i_b(w_sum_631), .i_c(w_sum_632), .ow_sum(w_sum_738), .ow_carry(w_carry_738));
wire w_sum_739, w_carry_739;
math_adder_carry_save CSA_739(.i_a(w_sum_476), .i_b(w_sum_477), .i_c(w_carry_631), .ow_sum(w_sum_739), .ow_carry(w_carry_739));
wire w_sum_740, w_carry_740;
math_adder_carry_save CSA_740(.i_a(w_carry_632), .i_b(w_sum_633), .i_c(w_sum_634), .ow_sum(w_sum_740), .ow_carry(w_carry_740));
wire w_sum_741, w_carry_741;
math_adder_carry_save CSA_741(.i_a(w_sum_480), .i_b(w_sum_481), .i_c(w_carry_633), .ow_sum(w_sum_741), .ow_carry(w_carry_741));
wire w_sum_742, w_carry_742;
math_adder_carry_save CSA_742(.i_a(w_carry_634), .i_b(w_sum_635), .i_c(w_sum_636), .ow_sum(w_sum_742), .ow_carry(w_carry_742));
wire w_sum_743, w_carry_743;
math_adder_carry_save CSA_743(.i_a(w_sum_484), .i_b(w_sum_485), .i_c(w_carry_635), .ow_sum(w_sum_743), .ow_carry(w_carry_743));
wire w_sum_744, w_carry_744;
math_adder_carry_save CSA_744(.i_a(w_carry_636), .i_b(w_sum_637), .i_c(w_sum_638), .ow_sum(w_sum_744), .ow_carry(w_carry_744));
wire w_sum_745, w_carry_745;
math_adder_carry_save CSA_745(.i_a(w_sum_488), .i_b(w_sum_489), .i_c(w_carry_637), .ow_sum(w_sum_745), .ow_carry(w_carry_745));
wire w_sum_746, w_carry_746;
math_adder_carry_save CSA_746(.i_a(w_carry_638), .i_b(w_sum_639), .i_c(w_sum_640), .ow_sum(w_sum_746), .ow_carry(w_carry_746));
wire w_sum_747, w_carry_747;
math_adder_carry_save CSA_747(.i_a(w_sum_492), .i_b(w_sum_493), .i_c(w_carry_639), .ow_sum(w_sum_747), .ow_carry(w_carry_747));
wire w_sum_748, w_carry_748;
math_adder_carry_save CSA_748(.i_a(w_carry_640), .i_b(w_sum_641), .i_c(w_sum_642), .ow_sum(w_sum_748), .ow_carry(w_carry_748));
wire w_sum_749, w_carry_749;
math_adder_carry_save CSA_749(.i_a(w_sum_496), .i_b(w_sum_497), .i_c(w_carry_641), .ow_sum(w_sum_749), .ow_carry(w_carry_749));
wire w_sum_750, w_carry_750;
math_adder_carry_save CSA_750(.i_a(w_carry_642), .i_b(w_sum_643), .i_c(w_sum_644), .ow_sum(w_sum_750), .ow_carry(w_carry_750));
wire w_sum_751, w_carry_751;
math_adder_carry_save CSA_751(.i_a(w_sum_500), .i_b(w_sum_501), .i_c(w_carry_643), .ow_sum(w_sum_751), .ow_carry(w_carry_751));
wire w_sum_752, w_carry_752;
math_adder_carry_save CSA_752(.i_a(w_carry_644), .i_b(w_sum_645), .i_c(w_sum_646), .ow_sum(w_sum_752), .ow_carry(w_carry_752));
wire w_sum_753, w_carry_753;
math_adder_carry_save CSA_753(.i_a(w_sum_504), .i_b(w_sum_505), .i_c(w_carry_645), .ow_sum(w_sum_753), .ow_carry(w_carry_753));
wire w_sum_754, w_carry_754;
math_adder_carry_save CSA_754(.i_a(w_carry_646), .i_b(w_sum_647), .i_c(w_sum_648), .ow_sum(w_sum_754), .ow_carry(w_carry_754));
wire w_sum_755, w_carry_755;
math_adder_carry_save CSA_755(.i_a(w_sum_508), .i_b(w_sum_509), .i_c(w_carry_647), .ow_sum(w_sum_755), .ow_carry(w_carry_755));
wire w_sum_756, w_carry_756;
math_adder_carry_save CSA_756(.i_a(w_carry_648), .i_b(w_sum_649), .i_c(w_sum_650), .ow_sum(w_sum_756), .ow_carry(w_carry_756));
wire w_sum_757, w_carry_757;
math_adder_carry_save CSA_757(.i_a(w_sum_512), .i_b(w_sum_513), .i_c(w_carry_649), .ow_sum(w_sum_757), .ow_carry(w_carry_757));
wire w_sum_758, w_carry_758;
math_adder_carry_save CSA_758(.i_a(w_carry_650), .i_b(w_sum_651), .i_c(w_sum_652), .ow_sum(w_sum_758), .ow_carry(w_carry_758));
wire w_sum_759, w_carry_759;
math_adder_carry_save CSA_759(.i_a(w_sum_516), .i_b(w_sum_517), .i_c(w_carry_651), .ow_sum(w_sum_759), .ow_carry(w_carry_759));
wire w_sum_760, w_carry_760;
math_adder_carry_save CSA_760(.i_a(w_carry_652), .i_b(w_sum_653), .i_c(w_sum_654), .ow_sum(w_sum_760), .ow_carry(w_carry_760));
wire w_sum_761, w_carry_761;
math_adder_carry_save CSA_761(.i_a(w_sum_520), .i_b(w_sum_521), .i_c(w_carry_653), .ow_sum(w_sum_761), .ow_carry(w_carry_761));
wire w_sum_762, w_carry_762;
math_adder_carry_save CSA_762(.i_a(w_carry_654), .i_b(w_sum_655), .i_c(w_sum_656), .ow_sum(w_sum_762), .ow_carry(w_carry_762));
wire w_sum_763, w_carry_763;
math_adder_carry_save CSA_763(.i_a(w_sum_524), .i_b(w_sum_525), .i_c(w_carry_655), .ow_sum(w_sum_763), .ow_carry(w_carry_763));
wire w_sum_764, w_carry_764;
math_adder_carry_save CSA_764(.i_a(w_carry_656), .i_b(w_sum_657), .i_c(w_sum_658), .ow_sum(w_sum_764), .ow_carry(w_carry_764));
wire w_sum_765, w_carry_765;
math_adder_carry_save CSA_765(.i_a(w_sum_528), .i_b(w_sum_529), .i_c(w_carry_657), .ow_sum(w_sum_765), .ow_carry(w_carry_765));
wire w_sum_766, w_carry_766;
math_adder_carry_save CSA_766(.i_a(w_carry_658), .i_b(w_sum_659), .i_c(w_sum_660), .ow_sum(w_sum_766), .ow_carry(w_carry_766));
wire w_sum_767, w_carry_767;
math_adder_carry_save CSA_767(.i_a(w_sum_532), .i_b(w_sum_533), .i_c(w_carry_659), .ow_sum(w_sum_767), .ow_carry(w_carry_767));
wire w_sum_768, w_carry_768;
math_adder_carry_save CSA_768(.i_a(w_carry_660), .i_b(w_sum_661), .i_c(w_sum_662), .ow_sum(w_sum_768), .ow_carry(w_carry_768));
wire w_sum_769, w_carry_769;
math_adder_carry_save CSA_769(.i_a(w_sum_536), .i_b(w_sum_537), .i_c(w_carry_661), .ow_sum(w_sum_769), .ow_carry(w_carry_769));
wire w_sum_770, w_carry_770;
math_adder_carry_save CSA_770(.i_a(w_carry_662), .i_b(w_sum_663), .i_c(w_sum_664), .ow_sum(w_sum_770), .ow_carry(w_carry_770));
wire w_sum_771, w_carry_771;
math_adder_carry_save CSA_771(.i_a(w_sum_540), .i_b(w_sum_541), .i_c(w_carry_663), .ow_sum(w_sum_771), .ow_carry(w_carry_771));
wire w_sum_772, w_carry_772;
math_adder_carry_save CSA_772(.i_a(w_carry_664), .i_b(w_sum_665), .i_c(w_sum_666), .ow_sum(w_sum_772), .ow_carry(w_carry_772));
wire w_sum_773, w_carry_773;
math_adder_carry_save CSA_773(.i_a(w_sum_544), .i_b(w_sum_545), .i_c(w_carry_665), .ow_sum(w_sum_773), .ow_carry(w_carry_773));
wire w_sum_774, w_carry_774;
math_adder_carry_save CSA_774(.i_a(w_carry_666), .i_b(w_sum_667), .i_c(w_sum_668), .ow_sum(w_sum_774), .ow_carry(w_carry_774));
wire w_sum_775, w_carry_775;
math_adder_carry_save CSA_775(.i_a(w_sum_548), .i_b(w_sum_549), .i_c(w_carry_667), .ow_sum(w_sum_775), .ow_carry(w_carry_775));
wire w_sum_776, w_carry_776;
math_adder_carry_save CSA_776(.i_a(w_carry_668), .i_b(w_sum_669), .i_c(w_sum_670), .ow_sum(w_sum_776), .ow_carry(w_carry_776));
wire w_sum_777, w_carry_777;
math_adder_carry_save CSA_777(.i_a(w_sum_552), .i_b(w_sum_553), .i_c(w_carry_669), .ow_sum(w_sum_777), .ow_carry(w_carry_777));
wire w_sum_778, w_carry_778;
math_adder_carry_save CSA_778(.i_a(w_carry_670), .i_b(w_sum_671), .i_c(w_sum_672), .ow_sum(w_sum_778), .ow_carry(w_carry_778));
wire w_sum_779, w_carry_779;
math_adder_carry_save CSA_779(.i_a(w_sum_556), .i_b(w_sum_557), .i_c(w_carry_671), .ow_sum(w_sum_779), .ow_carry(w_carry_779));
wire w_sum_780, w_carry_780;
math_adder_carry_save CSA_780(.i_a(w_carry_672), .i_b(w_sum_673), .i_c(w_sum_674), .ow_sum(w_sum_780), .ow_carry(w_carry_780));
wire w_sum_781, w_carry_781;
math_adder_carry_save CSA_781(.i_a(w_sum_560), .i_b(w_sum_561), .i_c(w_carry_673), .ow_sum(w_sum_781), .ow_carry(w_carry_781));
wire w_sum_782, w_carry_782;
math_adder_carry_save CSA_782(.i_a(w_carry_674), .i_b(w_sum_675), .i_c(w_sum_676), .ow_sum(w_sum_782), .ow_carry(w_carry_782));
wire w_sum_783, w_carry_783;
math_adder_carry_save CSA_783(.i_a(w_sum_564), .i_b(w_sum_565), .i_c(w_carry_675), .ow_sum(w_sum_783), .ow_carry(w_carry_783));
wire w_sum_784, w_carry_784;
math_adder_carry_save CSA_784(.i_a(w_carry_676), .i_b(w_sum_677), .i_c(w_sum_678), .ow_sum(w_sum_784), .ow_carry(w_carry_784));
wire w_sum_785, w_carry_785;
math_adder_carry_save CSA_785(.i_a(w_sum_568), .i_b(w_sum_569), .i_c(w_carry_677), .ow_sum(w_sum_785), .ow_carry(w_carry_785));
wire w_sum_786, w_carry_786;
math_adder_carry_save CSA_786(.i_a(w_carry_678), .i_b(w_sum_679), .i_c(w_sum_680), .ow_sum(w_sum_786), .ow_carry(w_carry_786));
wire w_sum_787, w_carry_787;
math_adder_carry_save CSA_787(.i_a(w_sum_572), .i_b(w_sum_573), .i_c(w_carry_679), .ow_sum(w_sum_787), .ow_carry(w_carry_787));
wire w_sum_788, w_carry_788;
math_adder_carry_save CSA_788(.i_a(w_carry_680), .i_b(w_sum_681), .i_c(w_sum_682), .ow_sum(w_sum_788), .ow_carry(w_carry_788));
wire w_sum_789, w_carry_789;
math_adder_carry_save CSA_789(.i_a(w_sum_576), .i_b(w_sum_577), .i_c(w_carry_681), .ow_sum(w_sum_789), .ow_carry(w_carry_789));
wire w_sum_790, w_carry_790;
math_adder_carry_save CSA_790(.i_a(w_carry_682), .i_b(w_sum_683), .i_c(w_sum_684), .ow_sum(w_sum_790), .ow_carry(w_carry_790));
wire w_sum_791, w_carry_791;
math_adder_carry_save CSA_791(.i_a(w_sum_580), .i_b(w_sum_581), .i_c(w_carry_683), .ow_sum(w_sum_791), .ow_carry(w_carry_791));
wire w_sum_792, w_carry_792;
math_adder_carry_save CSA_792(.i_a(w_carry_684), .i_b(w_sum_685), .i_c(w_sum_686), .ow_sum(w_sum_792), .ow_carry(w_carry_792));
wire w_sum_793, w_carry_793;
math_adder_carry_save CSA_793(.i_a(w_sum_584), .i_b(w_sum_585), .i_c(w_carry_685), .ow_sum(w_sum_793), .ow_carry(w_carry_793));
wire w_sum_794, w_carry_794;
math_adder_carry_save CSA_794(.i_a(w_carry_686), .i_b(w_sum_687), .i_c(w_sum_688), .ow_sum(w_sum_794), .ow_carry(w_carry_794));
wire w_sum_795, w_carry_795;
math_adder_carry_save CSA_795(.i_a(w_sum_588), .i_b(w_sum_589), .i_c(w_carry_687), .ow_sum(w_sum_795), .ow_carry(w_carry_795));
wire w_sum_796, w_carry_796;
math_adder_carry_save CSA_796(.i_a(w_carry_688), .i_b(w_sum_689), .i_c(w_sum_690), .ow_sum(w_sum_796), .ow_carry(w_carry_796));
wire w_sum_797, w_carry_797;
math_adder_carry_save CSA_797(.i_a(w_sum_592), .i_b(w_sum_593), .i_c(w_carry_689), .ow_sum(w_sum_797), .ow_carry(w_carry_797));
wire w_sum_798, w_carry_798;
math_adder_carry_save CSA_798(.i_a(w_carry_690), .i_b(w_sum_691), .i_c(w_sum_692), .ow_sum(w_sum_798), .ow_carry(w_carry_798));
wire w_sum_799, w_carry_799;
math_adder_carry_save CSA_799(.i_a(w_sum_595), .i_b(w_sum_596), .i_c(w_carry_691), .ow_sum(w_sum_799), .ow_carry(w_carry_799));
wire w_sum_800, w_carry_800;
math_adder_carry_save CSA_800(.i_a(w_carry_692), .i_b(w_sum_693), .i_c(w_sum_694), .ow_sum(w_sum_800), .ow_carry(w_carry_800));
wire w_sum_801, w_carry_801;
math_adder_carry_save CSA_801(.i_a(w_sum_597), .i_b(w_sum_598), .i_c(w_carry_693), .ow_sum(w_sum_801), .ow_carry(w_carry_801));
wire w_sum_802, w_carry_802;
math_adder_carry_save CSA_802(.i_a(w_carry_694), .i_b(w_sum_695), .i_c(w_sum_696), .ow_sum(w_sum_802), .ow_carry(w_carry_802));
wire w_sum_803, w_carry_803;
math_adder_carry_save CSA_803(.i_a(w_carry_598), .i_b(w_sum_599), .i_c(w_carry_695), .ow_sum(w_sum_803), .ow_carry(w_carry_803));
wire w_sum_804, w_carry_804;
math_adder_carry_save CSA_804(.i_a(w_carry_696), .i_b(w_sum_697), .i_c(w_sum_698), .ow_sum(w_sum_804), .ow_carry(w_carry_804));
wire w_sum_805, w_carry_805;
math_adder_carry_save CSA_805(.i_a(w_pp_31_25), .i_b(w_carry_599), .i_c(w_carry_697), .ow_sum(w_sum_805), .ow_carry(w_carry_805));
wire w_sum_806, w_carry_806;
math_adder_carry_save CSA_806(.i_a(w_carry_698), .i_b(w_sum_699), .i_c(w_sum_700), .ow_sum(w_sum_806), .ow_carry(w_carry_806));
wire w_sum_807, w_carry_807;
math_adder_carry_save CSA_807(.i_a(w_pp_29_28), .i_b(w_pp_30_27), .i_c(w_pp_31_26), .ow_sum(w_sum_807), .ow_carry(w_carry_807));
wire w_sum_808, w_carry_808;
math_adder_carry_save CSA_808(.i_a(w_carry_699), .i_b(w_carry_700), .i_c(w_sum_701), .ow_sum(w_sum_808), .ow_carry(w_carry_808));
wire w_sum_809, w_carry_809;
math_adder_carry_save CSA_809(.i_a(w_pp_27_31), .i_b(w_pp_28_30), .i_c(w_pp_29_29), .ow_sum(w_sum_809), .ow_carry(w_carry_809));
wire w_sum_810, w_carry_810;
math_adder_carry_save CSA_810(.i_a(w_pp_30_28), .i_b(w_pp_31_27), .i_c(w_carry_701), .ow_sum(w_sum_810), .ow_carry(w_carry_810));
wire w_sum_811, w_carry_811;
math_adder_carry_save CSA_811(.i_a(w_pp_28_31), .i_b(w_pp_29_30), .i_c(w_pp_30_29), .ow_sum(w_sum_811), .ow_carry(w_carry_811));
// Stage: 6, Max Height: 3
wire w_sum_812, w_carry_812;
math_adder_half HA_812(.i_a(w_pp_00_03), .i_b(w_pp_01_02), .ow_sum(w_sum_812), .ow_carry(w_carry_812));
wire w_sum_813, w_carry_813;
math_adder_carry_save CSA_813(.i_a(w_pp_02_02), .i_b(w_pp_03_01), .i_c(w_pp_04_00), .ow_sum(w_sum_813), .ow_carry(w_carry_813));
wire w_sum_814, w_carry_814;
math_adder_carry_save CSA_814(.i_a(w_pp_05_00), .i_b(w_carry_702), .i_c(w_sum_703), .ow_sum(w_sum_814), .ow_carry(w_carry_814));
wire w_sum_815, w_carry_815;
math_adder_carry_save CSA_815(.i_a(w_carry_703), .i_b(w_carry_704), .i_c(w_sum_705), .ow_sum(w_sum_815), .ow_carry(w_carry_815));
wire w_sum_816, w_carry_816;
math_adder_carry_save CSA_816(.i_a(w_carry_705), .i_b(w_carry_706), .i_c(w_sum_707), .ow_sum(w_sum_816), .ow_carry(w_carry_816));
wire w_sum_817, w_carry_817;
math_adder_carry_save CSA_817(.i_a(w_carry_707), .i_b(w_carry_708), .i_c(w_sum_709), .ow_sum(w_sum_817), .ow_carry(w_carry_817));
wire w_sum_818, w_carry_818;
math_adder_carry_save CSA_818(.i_a(w_carry_709), .i_b(w_carry_710), .i_c(w_sum_711), .ow_sum(w_sum_818), .ow_carry(w_carry_818));
wire w_sum_819, w_carry_819;
math_adder_carry_save CSA_819(.i_a(w_carry_711), .i_b(w_carry_712), .i_c(w_sum_713), .ow_sum(w_sum_819), .ow_carry(w_carry_819));
wire w_sum_820, w_carry_820;
math_adder_carry_save CSA_820(.i_a(w_carry_713), .i_b(w_carry_714), .i_c(w_sum_715), .ow_sum(w_sum_820), .ow_carry(w_carry_820));
wire w_sum_821, w_carry_821;
math_adder_carry_save CSA_821(.i_a(w_carry_715), .i_b(w_carry_716), .i_c(w_sum_717), .ow_sum(w_sum_821), .ow_carry(w_carry_821));
wire w_sum_822, w_carry_822;
math_adder_carry_save CSA_822(.i_a(w_carry_717), .i_b(w_carry_718), .i_c(w_sum_719), .ow_sum(w_sum_822), .ow_carry(w_carry_822));
wire w_sum_823, w_carry_823;
math_adder_carry_save CSA_823(.i_a(w_carry_719), .i_b(w_carry_720), .i_c(w_sum_721), .ow_sum(w_sum_823), .ow_carry(w_carry_823));
wire w_sum_824, w_carry_824;
math_adder_carry_save CSA_824(.i_a(w_carry_721), .i_b(w_carry_722), .i_c(w_sum_723), .ow_sum(w_sum_824), .ow_carry(w_carry_824));
wire w_sum_825, w_carry_825;
math_adder_carry_save CSA_825(.i_a(w_carry_723), .i_b(w_carry_724), .i_c(w_sum_725), .ow_sum(w_sum_825), .ow_carry(w_carry_825));
wire w_sum_826, w_carry_826;
math_adder_carry_save CSA_826(.i_a(w_carry_725), .i_b(w_carry_726), .i_c(w_sum_727), .ow_sum(w_sum_826), .ow_carry(w_carry_826));
wire w_sum_827, w_carry_827;
math_adder_carry_save CSA_827(.i_a(w_carry_727), .i_b(w_carry_728), .i_c(w_sum_729), .ow_sum(w_sum_827), .ow_carry(w_carry_827));
wire w_sum_828, w_carry_828;
math_adder_carry_save CSA_828(.i_a(w_carry_729), .i_b(w_carry_730), .i_c(w_sum_731), .ow_sum(w_sum_828), .ow_carry(w_carry_828));
wire w_sum_829, w_carry_829;
math_adder_carry_save CSA_829(.i_a(w_carry_731), .i_b(w_carry_732), .i_c(w_sum_733), .ow_sum(w_sum_829), .ow_carry(w_carry_829));
wire w_sum_830, w_carry_830;
math_adder_carry_save CSA_830(.i_a(w_carry_733), .i_b(w_carry_734), .i_c(w_sum_735), .ow_sum(w_sum_830), .ow_carry(w_carry_830));
wire w_sum_831, w_carry_831;
math_adder_carry_save CSA_831(.i_a(w_carry_735), .i_b(w_carry_736), .i_c(w_sum_737), .ow_sum(w_sum_831), .ow_carry(w_carry_831));
wire w_sum_832, w_carry_832;
math_adder_carry_save CSA_832(.i_a(w_carry_737), .i_b(w_carry_738), .i_c(w_sum_739), .ow_sum(w_sum_832), .ow_carry(w_carry_832));
wire w_sum_833, w_carry_833;
math_adder_carry_save CSA_833(.i_a(w_carry_739), .i_b(w_carry_740), .i_c(w_sum_741), .ow_sum(w_sum_833), .ow_carry(w_carry_833));
wire w_sum_834, w_carry_834;
math_adder_carry_save CSA_834(.i_a(w_carry_741), .i_b(w_carry_742), .i_c(w_sum_743), .ow_sum(w_sum_834), .ow_carry(w_carry_834));
wire w_sum_835, w_carry_835;
math_adder_carry_save CSA_835(.i_a(w_carry_743), .i_b(w_carry_744), .i_c(w_sum_745), .ow_sum(w_sum_835), .ow_carry(w_carry_835));
wire w_sum_836, w_carry_836;
math_adder_carry_save CSA_836(.i_a(w_carry_745), .i_b(w_carry_746), .i_c(w_sum_747), .ow_sum(w_sum_836), .ow_carry(w_carry_836));
wire w_sum_837, w_carry_837;
math_adder_carry_save CSA_837(.i_a(w_carry_747), .i_b(w_carry_748), .i_c(w_sum_749), .ow_sum(w_sum_837), .ow_carry(w_carry_837));
wire w_sum_838, w_carry_838;
math_adder_carry_save CSA_838(.i_a(w_carry_749), .i_b(w_carry_750), .i_c(w_sum_751), .ow_sum(w_sum_838), .ow_carry(w_carry_838));
wire w_sum_839, w_carry_839;
math_adder_carry_save CSA_839(.i_a(w_carry_751), .i_b(w_carry_752), .i_c(w_sum_753), .ow_sum(w_sum_839), .ow_carry(w_carry_839));
wire w_sum_840, w_carry_840;
math_adder_carry_save CSA_840(.i_a(w_carry_753), .i_b(w_carry_754), .i_c(w_sum_755), .ow_sum(w_sum_840), .ow_carry(w_carry_840));
wire w_sum_841, w_carry_841;
math_adder_carry_save CSA_841(.i_a(w_carry_755), .i_b(w_carry_756), .i_c(w_sum_757), .ow_sum(w_sum_841), .ow_carry(w_carry_841));
wire w_sum_842, w_carry_842;
math_adder_carry_save CSA_842(.i_a(w_carry_757), .i_b(w_carry_758), .i_c(w_sum_759), .ow_sum(w_sum_842), .ow_carry(w_carry_842));
wire w_sum_843, w_carry_843;
math_adder_carry_save CSA_843(.i_a(w_carry_759), .i_b(w_carry_760), .i_c(w_sum_761), .ow_sum(w_sum_843), .ow_carry(w_carry_843));
wire w_sum_844, w_carry_844;
math_adder_carry_save CSA_844(.i_a(w_carry_761), .i_b(w_carry_762), .i_c(w_sum_763), .ow_sum(w_sum_844), .ow_carry(w_carry_844));
wire w_sum_845, w_carry_845;
math_adder_carry_save CSA_845(.i_a(w_carry_763), .i_b(w_carry_764), .i_c(w_sum_765), .ow_sum(w_sum_845), .ow_carry(w_carry_845));
wire w_sum_846, w_carry_846;
math_adder_carry_save CSA_846(.i_a(w_carry_765), .i_b(w_carry_766), .i_c(w_sum_767), .ow_sum(w_sum_846), .ow_carry(w_carry_846));
wire w_sum_847, w_carry_847;
math_adder_carry_save CSA_847(.i_a(w_carry_767), .i_b(w_carry_768), .i_c(w_sum_769), .ow_sum(w_sum_847), .ow_carry(w_carry_847));
wire w_sum_848, w_carry_848;
math_adder_carry_save CSA_848(.i_a(w_carry_769), .i_b(w_carry_770), .i_c(w_sum_771), .ow_sum(w_sum_848), .ow_carry(w_carry_848));
wire w_sum_849, w_carry_849;
math_adder_carry_save CSA_849(.i_a(w_carry_771), .i_b(w_carry_772), .i_c(w_sum_773), .ow_sum(w_sum_849), .ow_carry(w_carry_849));
wire w_sum_850, w_carry_850;
math_adder_carry_save CSA_850(.i_a(w_carry_773), .i_b(w_carry_774), .i_c(w_sum_775), .ow_sum(w_sum_850), .ow_carry(w_carry_850));
wire w_sum_851, w_carry_851;
math_adder_carry_save CSA_851(.i_a(w_carry_775), .i_b(w_carry_776), .i_c(w_sum_777), .ow_sum(w_sum_851), .ow_carry(w_carry_851));
wire w_sum_852, w_carry_852;
math_adder_carry_save CSA_852(.i_a(w_carry_777), .i_b(w_carry_778), .i_c(w_sum_779), .ow_sum(w_sum_852), .ow_carry(w_carry_852));
wire w_sum_853, w_carry_853;
math_adder_carry_save CSA_853(.i_a(w_carry_779), .i_b(w_carry_780), .i_c(w_sum_781), .ow_sum(w_sum_853), .ow_carry(w_carry_853));
wire w_sum_854, w_carry_854;
math_adder_carry_save CSA_854(.i_a(w_carry_781), .i_b(w_carry_782), .i_c(w_sum_783), .ow_sum(w_sum_854), .ow_carry(w_carry_854));
wire w_sum_855, w_carry_855;
math_adder_carry_save CSA_855(.i_a(w_carry_783), .i_b(w_carry_784), .i_c(w_sum_785), .ow_sum(w_sum_855), .ow_carry(w_carry_855));
wire w_sum_856, w_carry_856;
math_adder_carry_save CSA_856(.i_a(w_carry_785), .i_b(w_carry_786), .i_c(w_sum_787), .ow_sum(w_sum_856), .ow_carry(w_carry_856));
wire w_sum_857, w_carry_857;
math_adder_carry_save CSA_857(.i_a(w_carry_787), .i_b(w_carry_788), .i_c(w_sum_789), .ow_sum(w_sum_857), .ow_carry(w_carry_857));
wire w_sum_858, w_carry_858;
math_adder_carry_save CSA_858(.i_a(w_carry_789), .i_b(w_carry_790), .i_c(w_sum_791), .ow_sum(w_sum_858), .ow_carry(w_carry_858));
wire w_sum_859, w_carry_859;
math_adder_carry_save CSA_859(.i_a(w_carry_791), .i_b(w_carry_792), .i_c(w_sum_793), .ow_sum(w_sum_859), .ow_carry(w_carry_859));
wire w_sum_860, w_carry_860;
math_adder_carry_save CSA_860(.i_a(w_carry_793), .i_b(w_carry_794), .i_c(w_sum_795), .ow_sum(w_sum_860), .ow_carry(w_carry_860));
wire w_sum_861, w_carry_861;
math_adder_carry_save CSA_861(.i_a(w_carry_795), .i_b(w_carry_796), .i_c(w_sum_797), .ow_sum(w_sum_861), .ow_carry(w_carry_861));
wire w_sum_862, w_carry_862;
math_adder_carry_save CSA_862(.i_a(w_carry_797), .i_b(w_carry_798), .i_c(w_sum_799), .ow_sum(w_sum_862), .ow_carry(w_carry_862));
wire w_sum_863, w_carry_863;
math_adder_carry_save CSA_863(.i_a(w_carry_799), .i_b(w_carry_800), .i_c(w_sum_801), .ow_sum(w_sum_863), .ow_carry(w_carry_863));
wire w_sum_864, w_carry_864;
math_adder_carry_save CSA_864(.i_a(w_carry_801), .i_b(w_carry_802), .i_c(w_sum_803), .ow_sum(w_sum_864), .ow_carry(w_carry_864));
wire w_sum_865, w_carry_865;
math_adder_carry_save CSA_865(.i_a(w_carry_803), .i_b(w_carry_804), .i_c(w_sum_805), .ow_sum(w_sum_865), .ow_carry(w_carry_865));
wire w_sum_866, w_carry_866;
math_adder_carry_save CSA_866(.i_a(w_carry_805), .i_b(w_carry_806), .i_c(w_sum_807), .ow_sum(w_sum_866), .ow_carry(w_carry_866));
wire w_sum_867, w_carry_867;
math_adder_carry_save CSA_867(.i_a(w_carry_807), .i_b(w_carry_808), .i_c(w_sum_809), .ow_sum(w_sum_867), .ow_carry(w_carry_867));
wire w_sum_868, w_carry_868;
math_adder_carry_save CSA_868(.i_a(w_pp_31_28), .i_b(w_carry_809), .i_c(w_carry_810), .ow_sum(w_sum_868), .ow_carry(w_carry_868));
wire w_sum_869, w_carry_869;
math_adder_carry_save CSA_869(.i_a(w_pp_29_31), .i_b(w_pp_30_30), .i_c(w_pp_31_29), .ow_sum(w_sum_869), .ow_carry(w_carry_869));
// Stage: 7, Max Height: 2
wire w_sum_870, w_carry_870;
math_adder_half HA_870(.i_a(w_pp_00_02), .i_b(w_pp_01_01), .ow_sum(w_sum_870), .ow_carry(w_carry_870));
wire w_sum_871, w_carry_871;
math_adder_carry_save CSA_871(.i_a(w_pp_02_01), .i_b(w_pp_03_00), .i_c(w_sum_812), .ow_sum(w_sum_871), .ow_carry(w_carry_871));
wire w_sum_872, w_carry_872;
math_adder_carry_save CSA_872(.i_a(w_sum_702), .i_b(w_carry_812), .i_c(w_sum_813), .ow_sum(w_sum_872), .ow_carry(w_carry_872));
wire w_sum_873, w_carry_873;
math_adder_carry_save CSA_873(.i_a(w_sum_704), .i_b(w_carry_813), .i_c(w_sum_814), .ow_sum(w_sum_873), .ow_carry(w_carry_873));
wire w_sum_874, w_carry_874;
math_adder_carry_save CSA_874(.i_a(w_sum_706), .i_b(w_carry_814), .i_c(w_sum_815), .ow_sum(w_sum_874), .ow_carry(w_carry_874));
wire w_sum_875, w_carry_875;
math_adder_carry_save CSA_875(.i_a(w_sum_708), .i_b(w_carry_815), .i_c(w_sum_816), .ow_sum(w_sum_875), .ow_carry(w_carry_875));
wire w_sum_876, w_carry_876;
math_adder_carry_save CSA_876(.i_a(w_sum_710), .i_b(w_carry_816), .i_c(w_sum_817), .ow_sum(w_sum_876), .ow_carry(w_carry_876));
wire w_sum_877, w_carry_877;
math_adder_carry_save CSA_877(.i_a(w_sum_712), .i_b(w_carry_817), .i_c(w_sum_818), .ow_sum(w_sum_877), .ow_carry(w_carry_877));
wire w_sum_878, w_carry_878;
math_adder_carry_save CSA_878(.i_a(w_sum_714), .i_b(w_carry_818), .i_c(w_sum_819), .ow_sum(w_sum_878), .ow_carry(w_carry_878));
wire w_sum_879, w_carry_879;
math_adder_carry_save CSA_879(.i_a(w_sum_716), .i_b(w_carry_819), .i_c(w_sum_820), .ow_sum(w_sum_879), .ow_carry(w_carry_879));
wire w_sum_880, w_carry_880;
math_adder_carry_save CSA_880(.i_a(w_sum_718), .i_b(w_carry_820), .i_c(w_sum_821), .ow_sum(w_sum_880), .ow_carry(w_carry_880));
wire w_sum_881, w_carry_881;
math_adder_carry_save CSA_881(.i_a(w_sum_720), .i_b(w_carry_821), .i_c(w_sum_822), .ow_sum(w_sum_881), .ow_carry(w_carry_881));
wire w_sum_882, w_carry_882;
math_adder_carry_save CSA_882(.i_a(w_sum_722), .i_b(w_carry_822), .i_c(w_sum_823), .ow_sum(w_sum_882), .ow_carry(w_carry_882));
wire w_sum_883, w_carry_883;
math_adder_carry_save CSA_883(.i_a(w_sum_724), .i_b(w_carry_823), .i_c(w_sum_824), .ow_sum(w_sum_883), .ow_carry(w_carry_883));
wire w_sum_884, w_carry_884;
math_adder_carry_save CSA_884(.i_a(w_sum_726), .i_b(w_carry_824), .i_c(w_sum_825), .ow_sum(w_sum_884), .ow_carry(w_carry_884));
wire w_sum_885, w_carry_885;
math_adder_carry_save CSA_885(.i_a(w_sum_728), .i_b(w_carry_825), .i_c(w_sum_826), .ow_sum(w_sum_885), .ow_carry(w_carry_885));
wire w_sum_886, w_carry_886;
math_adder_carry_save CSA_886(.i_a(w_sum_730), .i_b(w_carry_826), .i_c(w_sum_827), .ow_sum(w_sum_886), .ow_carry(w_carry_886));
wire w_sum_887, w_carry_887;
math_adder_carry_save CSA_887(.i_a(w_sum_732), .i_b(w_carry_827), .i_c(w_sum_828), .ow_sum(w_sum_887), .ow_carry(w_carry_887));
wire w_sum_888, w_carry_888;
math_adder_carry_save CSA_888(.i_a(w_sum_734), .i_b(w_carry_828), .i_c(w_sum_829), .ow_sum(w_sum_888), .ow_carry(w_carry_888));
wire w_sum_889, w_carry_889;
math_adder_carry_save CSA_889(.i_a(w_sum_736), .i_b(w_carry_829), .i_c(w_sum_830), .ow_sum(w_sum_889), .ow_carry(w_carry_889));
wire w_sum_890, w_carry_890;
math_adder_carry_save CSA_890(.i_a(w_sum_738), .i_b(w_carry_830), .i_c(w_sum_831), .ow_sum(w_sum_890), .ow_carry(w_carry_890));
wire w_sum_891, w_carry_891;
math_adder_carry_save CSA_891(.i_a(w_sum_740), .i_b(w_carry_831), .i_c(w_sum_832), .ow_sum(w_sum_891), .ow_carry(w_carry_891));
wire w_sum_892, w_carry_892;
math_adder_carry_save CSA_892(.i_a(w_sum_742), .i_b(w_carry_832), .i_c(w_sum_833), .ow_sum(w_sum_892), .ow_carry(w_carry_892));
wire w_sum_893, w_carry_893;
math_adder_carry_save CSA_893(.i_a(w_sum_744), .i_b(w_carry_833), .i_c(w_sum_834), .ow_sum(w_sum_893), .ow_carry(w_carry_893));
wire w_sum_894, w_carry_894;
math_adder_carry_save CSA_894(.i_a(w_sum_746), .i_b(w_carry_834), .i_c(w_sum_835), .ow_sum(w_sum_894), .ow_carry(w_carry_894));
wire w_sum_895, w_carry_895;
math_adder_carry_save CSA_895(.i_a(w_sum_748), .i_b(w_carry_835), .i_c(w_sum_836), .ow_sum(w_sum_895), .ow_carry(w_carry_895));
wire w_sum_896, w_carry_896;
math_adder_carry_save CSA_896(.i_a(w_sum_750), .i_b(w_carry_836), .i_c(w_sum_837), .ow_sum(w_sum_896), .ow_carry(w_carry_896));
wire w_sum_897, w_carry_897;
math_adder_carry_save CSA_897(.i_a(w_sum_752), .i_b(w_carry_837), .i_c(w_sum_838), .ow_sum(w_sum_897), .ow_carry(w_carry_897));
wire w_sum_898, w_carry_898;
math_adder_carry_save CSA_898(.i_a(w_sum_754), .i_b(w_carry_838), .i_c(w_sum_839), .ow_sum(w_sum_898), .ow_carry(w_carry_898));
wire w_sum_899, w_carry_899;
math_adder_carry_save CSA_899(.i_a(w_sum_756), .i_b(w_carry_839), .i_c(w_sum_840), .ow_sum(w_sum_899), .ow_carry(w_carry_899));
wire w_sum_900, w_carry_900;
math_adder_carry_save CSA_900(.i_a(w_sum_758), .i_b(w_carry_840), .i_c(w_sum_841), .ow_sum(w_sum_900), .ow_carry(w_carry_900));
wire w_sum_901, w_carry_901;
math_adder_carry_save CSA_901(.i_a(w_sum_760), .i_b(w_carry_841), .i_c(w_sum_842), .ow_sum(w_sum_901), .ow_carry(w_carry_901));
wire w_sum_902, w_carry_902;
math_adder_carry_save CSA_902(.i_a(w_sum_762), .i_b(w_carry_842), .i_c(w_sum_843), .ow_sum(w_sum_902), .ow_carry(w_carry_902));
wire w_sum_903, w_carry_903;
math_adder_carry_save CSA_903(.i_a(w_sum_764), .i_b(w_carry_843), .i_c(w_sum_844), .ow_sum(w_sum_903), .ow_carry(w_carry_903));
wire w_sum_904, w_carry_904;
math_adder_carry_save CSA_904(.i_a(w_sum_766), .i_b(w_carry_844), .i_c(w_sum_845), .ow_sum(w_sum_904), .ow_carry(w_carry_904));
wire w_sum_905, w_carry_905;
math_adder_carry_save CSA_905(.i_a(w_sum_768), .i_b(w_carry_845), .i_c(w_sum_846), .ow_sum(w_sum_905), .ow_carry(w_carry_905));
wire w_sum_906, w_carry_906;
math_adder_carry_save CSA_906(.i_a(w_sum_770), .i_b(w_carry_846), .i_c(w_sum_847), .ow_sum(w_sum_906), .ow_carry(w_carry_906));
wire w_sum_907, w_carry_907;
math_adder_carry_save CSA_907(.i_a(w_sum_772), .i_b(w_carry_847), .i_c(w_sum_848), .ow_sum(w_sum_907), .ow_carry(w_carry_907));
wire w_sum_908, w_carry_908;
math_adder_carry_save CSA_908(.i_a(w_sum_774), .i_b(w_carry_848), .i_c(w_sum_849), .ow_sum(w_sum_908), .ow_carry(w_carry_908));
wire w_sum_909, w_carry_909;
math_adder_carry_save CSA_909(.i_a(w_sum_776), .i_b(w_carry_849), .i_c(w_sum_850), .ow_sum(w_sum_909), .ow_carry(w_carry_909));
wire w_sum_910, w_carry_910;
math_adder_carry_save CSA_910(.i_a(w_sum_778), .i_b(w_carry_850), .i_c(w_sum_851), .ow_sum(w_sum_910), .ow_carry(w_carry_910));
wire w_sum_911, w_carry_911;
math_adder_carry_save CSA_911(.i_a(w_sum_780), .i_b(w_carry_851), .i_c(w_sum_852), .ow_sum(w_sum_911), .ow_carry(w_carry_911));
wire w_sum_912, w_carry_912;
math_adder_carry_save CSA_912(.i_a(w_sum_782), .i_b(w_carry_852), .i_c(w_sum_853), .ow_sum(w_sum_912), .ow_carry(w_carry_912));
wire w_sum_913, w_carry_913;
math_adder_carry_save CSA_913(.i_a(w_sum_784), .i_b(w_carry_853), .i_c(w_sum_854), .ow_sum(w_sum_913), .ow_carry(w_carry_913));
wire w_sum_914, w_carry_914;
math_adder_carry_save CSA_914(.i_a(w_sum_786), .i_b(w_carry_854), .i_c(w_sum_855), .ow_sum(w_sum_914), .ow_carry(w_carry_914));
wire w_sum_915, w_carry_915;
math_adder_carry_save CSA_915(.i_a(w_sum_788), .i_b(w_carry_855), .i_c(w_sum_856), .ow_sum(w_sum_915), .ow_carry(w_carry_915));
wire w_sum_916, w_carry_916;
math_adder_carry_save CSA_916(.i_a(w_sum_790), .i_b(w_carry_856), .i_c(w_sum_857), .ow_sum(w_sum_916), .ow_carry(w_carry_916));
wire w_sum_917, w_carry_917;
math_adder_carry_save CSA_917(.i_a(w_sum_792), .i_b(w_carry_857), .i_c(w_sum_858), .ow_sum(w_sum_917), .ow_carry(w_carry_917));
wire w_sum_918, w_carry_918;
math_adder_carry_save CSA_918(.i_a(w_sum_794), .i_b(w_carry_858), .i_c(w_sum_859), .ow_sum(w_sum_918), .ow_carry(w_carry_918));
wire w_sum_919, w_carry_919;
math_adder_carry_save CSA_919(.i_a(w_sum_796), .i_b(w_carry_859), .i_c(w_sum_860), .ow_sum(w_sum_919), .ow_carry(w_carry_919));
wire w_sum_920, w_carry_920;
math_adder_carry_save CSA_920(.i_a(w_sum_798), .i_b(w_carry_860), .i_c(w_sum_861), .ow_sum(w_sum_920), .ow_carry(w_carry_920));
wire w_sum_921, w_carry_921;
math_adder_carry_save CSA_921(.i_a(w_sum_800), .i_b(w_carry_861), .i_c(w_sum_862), .ow_sum(w_sum_921), .ow_carry(w_carry_921));
wire w_sum_922, w_carry_922;
math_adder_carry_save CSA_922(.i_a(w_sum_802), .i_b(w_carry_862), .i_c(w_sum_863), .ow_sum(w_sum_922), .ow_carry(w_carry_922));
wire w_sum_923, w_carry_923;
math_adder_carry_save CSA_923(.i_a(w_sum_804), .i_b(w_carry_863), .i_c(w_sum_864), .ow_sum(w_sum_923), .ow_carry(w_carry_923));
wire w_sum_924, w_carry_924;
math_adder_carry_save CSA_924(.i_a(w_sum_806), .i_b(w_carry_864), .i_c(w_sum_865), .ow_sum(w_sum_924), .ow_carry(w_carry_924));
wire w_sum_925, w_carry_925;
math_adder_carry_save CSA_925(.i_a(w_sum_808), .i_b(w_carry_865), .i_c(w_sum_866), .ow_sum(w_sum_925), .ow_carry(w_carry_925));
wire w_sum_926, w_carry_926;
math_adder_carry_save CSA_926(.i_a(w_sum_810), .i_b(w_carry_866), .i_c(w_sum_867), .ow_sum(w_sum_926), .ow_carry(w_carry_926));
wire w_sum_927, w_carry_927;
math_adder_carry_save CSA_927(.i_a(w_sum_811), .i_b(w_carry_867), .i_c(w_sum_868), .ow_sum(w_sum_927), .ow_carry(w_carry_927));
wire w_sum_928, w_carry_928;
math_adder_carry_save CSA_928(.i_a(w_carry_811), .i_b(w_carry_868), .i_c(w_sum_869), .ow_sum(w_sum_928), .ow_carry(w_carry_928));
wire w_sum_929, w_carry_929;
math_adder_carry_save CSA_929(.i_a(w_pp_30_31), .i_b(w_pp_31_30), .i_c(w_carry_869), .ow_sum(w_sum_929), .ow_carry(w_carry_929));

// Final addition stage
wire ow_sum_00, ow_carry_00;
assign ow_sum_00 = w_pp_00_00;
assign ow_carry_00 = 1'b0;
wire ow_sum_01, ow_carry_01;
math_adder_full FA_01(.i_a(w_pp_00_01), .i_b(w_pp_01_00), .i_c(ow_carry_00), .ow_sum(ow_sum_01), .ow_carry(ow_carry_01));
wire ow_sum_02, ow_carry_02;
math_adder_full FA_02(.i_a(w_pp_02_00), .i_b(w_sum_870), .i_c(ow_carry_01), .ow_sum(ow_sum_02), .ow_carry(ow_carry_02));
wire ow_sum_03, ow_carry_03;
math_adder_full FA_03(.i_a(w_carry_870), .i_b(w_sum_871), .i_c(ow_carry_02), .ow_sum(ow_sum_03), .ow_carry(ow_carry_03));
wire ow_sum_04, ow_carry_04;
math_adder_full FA_04(.i_a(w_carry_871), .i_b(w_sum_872), .i_c(ow_carry_03), .ow_sum(ow_sum_04), .ow_carry(ow_carry_04));
wire ow_sum_05, ow_carry_05;
math_adder_full FA_05(.i_a(w_carry_872), .i_b(w_sum_873), .i_c(ow_carry_04), .ow_sum(ow_sum_05), .ow_carry(ow_carry_05));
wire ow_sum_06, ow_carry_06;
math_adder_full FA_06(.i_a(w_carry_873), .i_b(w_sum_874), .i_c(ow_carry_05), .ow_sum(ow_sum_06), .ow_carry(ow_carry_06));
wire ow_sum_07, ow_carry_07;
math_adder_full FA_07(.i_a(w_carry_874), .i_b(w_sum_875), .i_c(ow_carry_06), .ow_sum(ow_sum_07), .ow_carry(ow_carry_07));
wire ow_sum_08, ow_carry_08;
math_adder_full FA_08(.i_a(w_carry_875), .i_b(w_sum_876), .i_c(ow_carry_07), .ow_sum(ow_sum_08), .ow_carry(ow_carry_08));
wire ow_sum_09, ow_carry_09;
math_adder_full FA_09(.i_a(w_carry_876), .i_b(w_sum_877), .i_c(ow_carry_08), .ow_sum(ow_sum_09), .ow_carry(ow_carry_09));
wire ow_sum_10, ow_carry_10;
math_adder_full FA_10(.i_a(w_carry_877), .i_b(w_sum_878), .i_c(ow_carry_09), .ow_sum(ow_sum_10), .ow_carry(ow_carry_10));
wire ow_sum_11, ow_carry_11;
math_adder_full FA_11(.i_a(w_carry_878), .i_b(w_sum_879), .i_c(ow_carry_10), .ow_sum(ow_sum_11), .ow_carry(ow_carry_11));
wire ow_sum_12, ow_carry_12;
math_adder_full FA_12(.i_a(w_carry_879), .i_b(w_sum_880), .i_c(ow_carry_11), .ow_sum(ow_sum_12), .ow_carry(ow_carry_12));
wire ow_sum_13, ow_carry_13;
math_adder_full FA_13(.i_a(w_carry_880), .i_b(w_sum_881), .i_c(ow_carry_12), .ow_sum(ow_sum_13), .ow_carry(ow_carry_13));
wire ow_sum_14, ow_carry_14;
math_adder_full FA_14(.i_a(w_carry_881), .i_b(w_sum_882), .i_c(ow_carry_13), .ow_sum(ow_sum_14), .ow_carry(ow_carry_14));
wire ow_sum_15, ow_carry_15;
math_adder_full FA_15(.i_a(w_carry_882), .i_b(w_sum_883), .i_c(ow_carry_14), .ow_sum(ow_sum_15), .ow_carry(ow_carry_15));
wire ow_sum_16, ow_carry_16;
math_adder_full FA_16(.i_a(w_carry_883), .i_b(w_sum_884), .i_c(ow_carry_15), .ow_sum(ow_sum_16), .ow_carry(ow_carry_16));
wire ow_sum_17, ow_carry_17;
math_adder_full FA_17(.i_a(w_carry_884), .i_b(w_sum_885), .i_c(ow_carry_16), .ow_sum(ow_sum_17), .ow_carry(ow_carry_17));
wire ow_sum_18, ow_carry_18;
math_adder_full FA_18(.i_a(w_carry_885), .i_b(w_sum_886), .i_c(ow_carry_17), .ow_sum(ow_sum_18), .ow_carry(ow_carry_18));
wire ow_sum_19, ow_carry_19;
math_adder_full FA_19(.i_a(w_carry_886), .i_b(w_sum_887), .i_c(ow_carry_18), .ow_sum(ow_sum_19), .ow_carry(ow_carry_19));
wire ow_sum_20, ow_carry_20;
math_adder_full FA_20(.i_a(w_carry_887), .i_b(w_sum_888), .i_c(ow_carry_19), .ow_sum(ow_sum_20), .ow_carry(ow_carry_20));
wire ow_sum_21, ow_carry_21;
math_adder_full FA_21(.i_a(w_carry_888), .i_b(w_sum_889), .i_c(ow_carry_20), .ow_sum(ow_sum_21), .ow_carry(ow_carry_21));
wire ow_sum_22, ow_carry_22;
math_adder_full FA_22(.i_a(w_carry_889), .i_b(w_sum_890), .i_c(ow_carry_21), .ow_sum(ow_sum_22), .ow_carry(ow_carry_22));
wire ow_sum_23, ow_carry_23;
math_adder_full FA_23(.i_a(w_carry_890), .i_b(w_sum_891), .i_c(ow_carry_22), .ow_sum(ow_sum_23), .ow_carry(ow_carry_23));
wire ow_sum_24, ow_carry_24;
math_adder_full FA_24(.i_a(w_carry_891), .i_b(w_sum_892), .i_c(ow_carry_23), .ow_sum(ow_sum_24), .ow_carry(ow_carry_24));
wire ow_sum_25, ow_carry_25;
math_adder_full FA_25(.i_a(w_carry_892), .i_b(w_sum_893), .i_c(ow_carry_24), .ow_sum(ow_sum_25), .ow_carry(ow_carry_25));
wire ow_sum_26, ow_carry_26;
math_adder_full FA_26(.i_a(w_carry_893), .i_b(w_sum_894), .i_c(ow_carry_25), .ow_sum(ow_sum_26), .ow_carry(ow_carry_26));
wire ow_sum_27, ow_carry_27;
math_adder_full FA_27(.i_a(w_carry_894), .i_b(w_sum_895), .i_c(ow_carry_26), .ow_sum(ow_sum_27), .ow_carry(ow_carry_27));
wire ow_sum_28, ow_carry_28;
math_adder_full FA_28(.i_a(w_carry_895), .i_b(w_sum_896), .i_c(ow_carry_27), .ow_sum(ow_sum_28), .ow_carry(ow_carry_28));
wire ow_sum_29, ow_carry_29;
math_adder_full FA_29(.i_a(w_carry_896), .i_b(w_sum_897), .i_c(ow_carry_28), .ow_sum(ow_sum_29), .ow_carry(ow_carry_29));
wire ow_sum_30, ow_carry_30;
math_adder_full FA_30(.i_a(w_carry_897), .i_b(w_sum_898), .i_c(ow_carry_29), .ow_sum(ow_sum_30), .ow_carry(ow_carry_30));
wire ow_sum_31, ow_carry_31;
math_adder_full FA_31(.i_a(w_carry_898), .i_b(w_sum_899), .i_c(ow_carry_30), .ow_sum(ow_sum_31), .ow_carry(ow_carry_31));
wire ow_sum_32, ow_carry_32;
math_adder_full FA_32(.i_a(w_carry_899), .i_b(w_sum_900), .i_c(ow_carry_31), .ow_sum(ow_sum_32), .ow_carry(ow_carry_32));
wire ow_sum_33, ow_carry_33;
math_adder_full FA_33(.i_a(w_carry_900), .i_b(w_sum_901), .i_c(ow_carry_32), .ow_sum(ow_sum_33), .ow_carry(ow_carry_33));
wire ow_sum_34, ow_carry_34;
math_adder_full FA_34(.i_a(w_carry_901), .i_b(w_sum_902), .i_c(ow_carry_33), .ow_sum(ow_sum_34), .ow_carry(ow_carry_34));
wire ow_sum_35, ow_carry_35;
math_adder_full FA_35(.i_a(w_carry_902), .i_b(w_sum_903), .i_c(ow_carry_34), .ow_sum(ow_sum_35), .ow_carry(ow_carry_35));
wire ow_sum_36, ow_carry_36;
math_adder_full FA_36(.i_a(w_carry_903), .i_b(w_sum_904), .i_c(ow_carry_35), .ow_sum(ow_sum_36), .ow_carry(ow_carry_36));
wire ow_sum_37, ow_carry_37;
math_adder_full FA_37(.i_a(w_carry_904), .i_b(w_sum_905), .i_c(ow_carry_36), .ow_sum(ow_sum_37), .ow_carry(ow_carry_37));
wire ow_sum_38, ow_carry_38;
math_adder_full FA_38(.i_a(w_carry_905), .i_b(w_sum_906), .i_c(ow_carry_37), .ow_sum(ow_sum_38), .ow_carry(ow_carry_38));
wire ow_sum_39, ow_carry_39;
math_adder_full FA_39(.i_a(w_carry_906), .i_b(w_sum_907), .i_c(ow_carry_38), .ow_sum(ow_sum_39), .ow_carry(ow_carry_39));
wire ow_sum_40, ow_carry_40;
math_adder_full FA_40(.i_a(w_carry_907), .i_b(w_sum_908), .i_c(ow_carry_39), .ow_sum(ow_sum_40), .ow_carry(ow_carry_40));
wire ow_sum_41, ow_carry_41;
math_adder_full FA_41(.i_a(w_carry_908), .i_b(w_sum_909), .i_c(ow_carry_40), .ow_sum(ow_sum_41), .ow_carry(ow_carry_41));
wire ow_sum_42, ow_carry_42;
math_adder_full FA_42(.i_a(w_carry_909), .i_b(w_sum_910), .i_c(ow_carry_41), .ow_sum(ow_sum_42), .ow_carry(ow_carry_42));
wire ow_sum_43, ow_carry_43;
math_adder_full FA_43(.i_a(w_carry_910), .i_b(w_sum_911), .i_c(ow_carry_42), .ow_sum(ow_sum_43), .ow_carry(ow_carry_43));
wire ow_sum_44, ow_carry_44;
math_adder_full FA_44(.i_a(w_carry_911), .i_b(w_sum_912), .i_c(ow_carry_43), .ow_sum(ow_sum_44), .ow_carry(ow_carry_44));
wire ow_sum_45, ow_carry_45;
math_adder_full FA_45(.i_a(w_carry_912), .i_b(w_sum_913), .i_c(ow_carry_44), .ow_sum(ow_sum_45), .ow_carry(ow_carry_45));
wire ow_sum_46, ow_carry_46;
math_adder_full FA_46(.i_a(w_carry_913), .i_b(w_sum_914), .i_c(ow_carry_45), .ow_sum(ow_sum_46), .ow_carry(ow_carry_46));
wire ow_sum_47, ow_carry_47;
math_adder_full FA_47(.i_a(w_carry_914), .i_b(w_sum_915), .i_c(ow_carry_46), .ow_sum(ow_sum_47), .ow_carry(ow_carry_47));
wire ow_sum_48, ow_carry_48;
math_adder_full FA_48(.i_a(w_carry_915), .i_b(w_sum_916), .i_c(ow_carry_47), .ow_sum(ow_sum_48), .ow_carry(ow_carry_48));
wire ow_sum_49, ow_carry_49;
math_adder_full FA_49(.i_a(w_carry_916), .i_b(w_sum_917), .i_c(ow_carry_48), .ow_sum(ow_sum_49), .ow_carry(ow_carry_49));
wire ow_sum_50, ow_carry_50;
math_adder_full FA_50(.i_a(w_carry_917), .i_b(w_sum_918), .i_c(ow_carry_49), .ow_sum(ow_sum_50), .ow_carry(ow_carry_50));
wire ow_sum_51, ow_carry_51;
math_adder_full FA_51(.i_a(w_carry_918), .i_b(w_sum_919), .i_c(ow_carry_50), .ow_sum(ow_sum_51), .ow_carry(ow_carry_51));
wire ow_sum_52, ow_carry_52;
math_adder_full FA_52(.i_a(w_carry_919), .i_b(w_sum_920), .i_c(ow_carry_51), .ow_sum(ow_sum_52), .ow_carry(ow_carry_52));
wire ow_sum_53, ow_carry_53;
math_adder_full FA_53(.i_a(w_carry_920), .i_b(w_sum_921), .i_c(ow_carry_52), .ow_sum(ow_sum_53), .ow_carry(ow_carry_53));
wire ow_sum_54, ow_carry_54;
math_adder_full FA_54(.i_a(w_carry_921), .i_b(w_sum_922), .i_c(ow_carry_53), .ow_sum(ow_sum_54), .ow_carry(ow_carry_54));
wire ow_sum_55, ow_carry_55;
math_adder_full FA_55(.i_a(w_carry_922), .i_b(w_sum_923), .i_c(ow_carry_54), .ow_sum(ow_sum_55), .ow_carry(ow_carry_55));
wire ow_sum_56, ow_carry_56;
math_adder_full FA_56(.i_a(w_carry_923), .i_b(w_sum_924), .i_c(ow_carry_55), .ow_sum(ow_sum_56), .ow_carry(ow_carry_56));
wire ow_sum_57, ow_carry_57;
math_adder_full FA_57(.i_a(w_carry_924), .i_b(w_sum_925), .i_c(ow_carry_56), .ow_sum(ow_sum_57), .ow_carry(ow_carry_57));
wire ow_sum_58, ow_carry_58;
math_adder_full FA_58(.i_a(w_carry_925), .i_b(w_sum_926), .i_c(ow_carry_57), .ow_sum(ow_sum_58), .ow_carry(ow_carry_58));
wire ow_sum_59, ow_carry_59;
math_adder_full FA_59(.i_a(w_carry_926), .i_b(w_sum_927), .i_c(ow_carry_58), .ow_sum(ow_sum_59), .ow_carry(ow_carry_59));
wire ow_sum_60, ow_carry_60;
math_adder_full FA_60(.i_a(w_carry_927), .i_b(w_sum_928), .i_c(ow_carry_59), .ow_sum(ow_sum_60), .ow_carry(ow_carry_60));
wire ow_sum_61, ow_carry_61;
math_adder_full FA_61(.i_a(w_carry_928), .i_b(w_sum_929), .i_c(ow_carry_60), .ow_sum(ow_sum_61), .ow_carry(ow_carry_61));
wire ow_sum_62, ow_carry_62;
math_adder_full FA_62(.i_a(w_pp_31_31), .i_b(w_carry_929), .i_c(ow_carry_61), .ow_sum(ow_sum_62), .ow_carry(ow_carry_62));
wire ow_sum_63, ow_carry_63;
assign ow_sum_63 = ow_carry_62;
assign ow_carry_63 = 1'b0;

// Final product assignment
assign ow_product[ 0] = ow_sum_00;
assign ow_product[ 1] = ow_sum_01;
assign ow_product[ 2] = ow_sum_02;
assign ow_product[ 3] = ow_sum_03;
assign ow_product[ 4] = ow_sum_04;
assign ow_product[ 5] = ow_sum_05;
assign ow_product[ 6] = ow_sum_06;
assign ow_product[ 7] = ow_sum_07;
assign ow_product[ 8] = ow_sum_08;
assign ow_product[ 9] = ow_sum_09;
assign ow_product[10] = ow_sum_10;
assign ow_product[11] = ow_sum_11;
assign ow_product[12] = ow_sum_12;
assign ow_product[13] = ow_sum_13;
assign ow_product[14] = ow_sum_14;
assign ow_product[15] = ow_sum_15;
assign ow_product[16] = ow_sum_16;
assign ow_product[17] = ow_sum_17;
assign ow_product[18] = ow_sum_18;
assign ow_product[19] = ow_sum_19;
assign ow_product[20] = ow_sum_20;
assign ow_product[21] = ow_sum_21;
assign ow_product[22] = ow_sum_22;
assign ow_product[23] = ow_sum_23;
assign ow_product[24] = ow_sum_24;
assign ow_product[25] = ow_sum_25;
assign ow_product[26] = ow_sum_26;
assign ow_product[27] = ow_sum_27;
assign ow_product[28] = ow_sum_28;
assign ow_product[29] = ow_sum_29;
assign ow_product[30] = ow_sum_30;
assign ow_product[31] = ow_sum_31;
assign ow_product[32] = ow_sum_32;
assign ow_product[33] = ow_sum_33;
assign ow_product[34] = ow_sum_34;
assign ow_product[35] = ow_sum_35;
assign ow_product[36] = ow_sum_36;
assign ow_product[37] = ow_sum_37;
assign ow_product[38] = ow_sum_38;
assign ow_product[39] = ow_sum_39;
assign ow_product[40] = ow_sum_40;
assign ow_product[41] = ow_sum_41;
assign ow_product[42] = ow_sum_42;
assign ow_product[43] = ow_sum_43;
assign ow_product[44] = ow_sum_44;
assign ow_product[45] = ow_sum_45;
assign ow_product[46] = ow_sum_46;
assign ow_product[47] = ow_sum_47;
assign ow_product[48] = ow_sum_48;
assign ow_product[49] = ow_sum_49;
assign ow_product[50] = ow_sum_50;
assign ow_product[51] = ow_sum_51;
assign ow_product[52] = ow_sum_52;
assign ow_product[53] = ow_sum_53;
assign ow_product[54] = ow_sum_54;
assign ow_product[55] = ow_sum_55;
assign ow_product[56] = ow_sum_56;
assign ow_product[57] = ow_sum_57;
assign ow_product[58] = ow_sum_58;
assign ow_product[59] = ow_sum_59;
assign ow_product[60] = ow_sum_60;
assign ow_product[61] = ow_sum_61;
assign ow_product[62] = ow_sum_62;
assign ow_product[63] = ow_sum_63;


    // Debug purposes
    // synopsys translate_off
    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, math_multiplier_dadda_tree_32);
    end
    // synopsys translate_off
        
endmodule : math_multiplier_dadda_tree_32
